VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fa16b_rev
  CLASS BLOCK ;
  FOREIGN 16b_FA ;
  ORIGIN 0.000 0.000 ;
  SIZE 150.000 BY 340.000 ;
  PIN c15_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 90.965 14.805 91.345 15.185 ;
        RECT 87.890 14.295 90.590 14.715 ;
        RECT 90.075 11.870 93.150 12.145 ;
        RECT 90.090 8.445 91.400 8.765 ;
        RECT 87.900 7.890 88.280 8.270 ;
      LAYER Metal2 ;
        RECT 87.940 7.800 88.240 14.740 ;
        RECT 90.150 8.375 90.455 14.735 ;
        RECT 91.000 8.375 91.300 15.195 ;
    END
  END c15_not
  PIN c15
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 84.065 14.815 84.445 15.195 ;
        RECT 81.390 14.390 83.130 14.680 ;
        RECT 82.745 9.795 93.150 10.130 ;
        RECT 82.715 8.475 84.495 8.765 ;
        RECT 81.445 7.860 81.825 8.240 ;
      LAYER Metal2 ;
        RECT 81.475 7.800 81.775 14.730 ;
        RECT 82.785 8.400 83.085 14.750 ;
        RECT 84.100 8.430 84.395 15.255 ;
    END
  END c15
  PIN s5_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 135.025 232.285 135.405 232.665 ;
        RECT 131.950 231.790 134.575 232.200 ;
        RECT 134.135 229.350 137.210 229.625 ;
        RECT 134.150 225.925 135.460 226.245 ;
        RECT 131.960 225.370 132.340 225.750 ;
      LAYER Metal2 ;
        RECT 132.000 225.280 132.300 232.220 ;
        RECT 134.210 225.855 134.490 232.215 ;
        RECT 135.060 225.855 135.360 232.675 ;
    END
  END s5_not
  PIN s5
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 128.125 232.295 128.505 232.675 ;
        RECT 125.450 231.870 127.190 232.160 ;
        RECT 126.805 227.275 137.210 227.610 ;
        RECT 126.775 225.955 128.555 226.245 ;
        RECT 125.505 225.340 125.885 225.720 ;
      LAYER Metal2 ;
        RECT 125.535 225.280 125.835 232.210 ;
        RECT 126.845 225.880 127.145 232.230 ;
        RECT 128.160 225.910 128.455 232.735 ;
    END
  END s5
  PIN s0_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 135.045 330.920 135.425 331.300 ;
        RECT 131.970 330.425 134.595 330.835 ;
        RECT 134.155 327.985 137.230 328.260 ;
        RECT 134.170 324.560 135.480 324.880 ;
        RECT 131.980 324.005 132.360 324.385 ;
      LAYER Metal2 ;
        RECT 132.020 323.915 132.320 330.855 ;
        RECT 134.230 324.490 134.510 330.850 ;
        RECT 135.080 324.490 135.380 331.310 ;
    END
  END s0_not
  PIN s0
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 128.145 330.930 128.525 331.310 ;
        RECT 125.470 330.505 127.210 330.795 ;
        RECT 126.825 325.910 137.230 326.245 ;
        RECT 126.795 324.590 128.575 324.880 ;
        RECT 125.525 323.975 125.905 324.355 ;
      LAYER Metal2 ;
        RECT 125.555 323.915 125.855 330.845 ;
        RECT 126.865 324.515 127.165 330.865 ;
        RECT 128.180 324.545 128.475 331.370 ;
    END
  END s0
  PIN s6_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 135.025 212.315 135.405 212.695 ;
        RECT 131.950 211.820 134.575 212.230 ;
        RECT 134.135 209.380 137.210 209.655 ;
        RECT 134.150 205.955 135.460 206.275 ;
        RECT 131.960 205.400 132.340 205.780 ;
      LAYER Metal2 ;
        RECT 132.000 205.310 132.300 212.250 ;
        RECT 134.210 205.885 134.490 212.245 ;
        RECT 135.060 205.885 135.360 212.705 ;
    END
  END s6_not
  PIN s6
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 128.125 212.325 128.505 212.705 ;
        RECT 125.450 211.900 127.190 212.190 ;
        RECT 126.805 207.305 137.210 207.640 ;
        RECT 126.775 205.985 128.555 206.275 ;
        RECT 125.505 205.370 125.885 205.750 ;
      LAYER Metal2 ;
        RECT 125.535 205.310 125.835 212.240 ;
        RECT 126.845 205.910 127.145 212.260 ;
        RECT 128.160 205.940 128.455 212.765 ;
    END
  END s6
  PIN s1_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 134.845 311.195 135.225 311.575 ;
        RECT 131.770 310.700 134.395 311.110 ;
        RECT 133.955 308.260 137.030 308.535 ;
        RECT 133.970 304.835 135.280 305.155 ;
        RECT 131.780 304.280 132.160 304.660 ;
      LAYER Metal2 ;
        RECT 131.820 304.190 132.120 311.130 ;
        RECT 134.030 304.765 134.310 311.125 ;
        RECT 134.880 304.765 135.180 311.585 ;
    END
  END s1_not
  PIN s1
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 127.945 311.205 128.325 311.585 ;
        RECT 125.270 310.780 127.010 311.070 ;
        RECT 126.625 306.185 137.030 306.520 ;
        RECT 126.595 304.865 128.375 305.155 ;
        RECT 125.325 304.250 125.705 304.630 ;
      LAYER Metal2 ;
        RECT 125.355 304.190 125.655 311.120 ;
        RECT 126.665 304.790 126.965 311.140 ;
        RECT 127.980 304.820 128.275 311.645 ;
    END
  END s1
  PIN s7_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 135.025 192.650 135.405 193.030 ;
        RECT 131.950 192.155 134.575 192.565 ;
        RECT 134.135 189.715 137.210 189.990 ;
        RECT 134.150 186.290 135.460 186.610 ;
        RECT 131.960 185.735 132.340 186.115 ;
      LAYER Metal2 ;
        RECT 132.000 185.645 132.300 192.585 ;
        RECT 134.210 186.220 134.490 192.580 ;
        RECT 135.060 186.220 135.360 193.040 ;
    END
  END s7_not
  PIN s7
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 128.125 192.660 128.505 193.040 ;
        RECT 125.450 192.235 127.190 192.525 ;
        RECT 126.805 187.640 137.210 187.975 ;
        RECT 126.775 186.320 128.555 186.610 ;
        RECT 125.505 185.705 125.885 186.085 ;
      LAYER Metal2 ;
        RECT 125.535 185.645 125.835 192.575 ;
        RECT 126.845 186.245 127.145 192.595 ;
        RECT 128.160 186.275 128.455 193.100 ;
    END
  END s7
  PIN s2_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 135.000 291.550 135.380 291.930 ;
        RECT 131.925 291.055 134.550 291.465 ;
        RECT 134.110 288.615 137.185 288.890 ;
        RECT 134.125 285.190 135.435 285.510 ;
        RECT 131.935 284.635 132.315 285.015 ;
      LAYER Metal2 ;
        RECT 131.975 284.545 132.275 291.485 ;
        RECT 134.185 285.120 134.465 291.480 ;
        RECT 135.035 285.120 135.335 291.940 ;
    END
  END s2_not
  PIN s2
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 128.100 291.560 128.480 291.940 ;
        RECT 125.425 291.135 127.165 291.425 ;
        RECT 126.780 286.540 137.185 286.875 ;
        RECT 126.750 285.220 128.530 285.510 ;
        RECT 125.480 284.605 125.860 284.985 ;
      LAYER Metal2 ;
        RECT 125.510 284.545 125.810 291.475 ;
        RECT 126.820 285.145 127.120 291.495 ;
        RECT 128.135 285.175 128.430 292.000 ;
    END
  END s2
  PIN s8_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 135.065 172.810 135.445 173.190 ;
        RECT 131.990 172.315 134.615 172.725 ;
        RECT 134.175 169.875 137.250 170.150 ;
        RECT 134.190 166.450 135.500 166.770 ;
        RECT 132.000 165.895 132.380 166.275 ;
      LAYER Metal2 ;
        RECT 132.040 165.805 132.340 172.745 ;
        RECT 134.250 166.380 134.530 172.740 ;
        RECT 135.100 166.380 135.400 173.200 ;
    END
  END s8_not
  PIN s8
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 128.165 172.820 128.545 173.200 ;
        RECT 125.490 172.395 127.230 172.685 ;
        RECT 126.845 167.800 137.250 168.135 ;
        RECT 126.815 166.480 128.595 166.770 ;
        RECT 125.545 165.865 125.925 166.245 ;
      LAYER Metal2 ;
        RECT 125.575 165.805 125.875 172.735 ;
        RECT 126.885 166.405 127.185 172.755 ;
        RECT 128.200 166.435 128.495 173.260 ;
    END
  END s8
  PIN s3_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 135.000 271.755 135.380 272.135 ;
        RECT 131.925 271.260 134.550 271.670 ;
        RECT 134.110 268.820 137.185 269.095 ;
        RECT 134.125 265.395 135.435 265.715 ;
        RECT 131.935 264.840 132.315 265.220 ;
      LAYER Metal2 ;
        RECT 131.975 264.750 132.275 271.690 ;
        RECT 134.185 265.325 134.465 271.685 ;
        RECT 135.035 265.325 135.335 272.145 ;
    END
  END s3_not
  PIN s3
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 128.100 271.765 128.480 272.145 ;
        RECT 125.425 271.340 127.165 271.630 ;
        RECT 126.780 266.745 137.185 267.080 ;
        RECT 126.750 265.425 128.530 265.715 ;
        RECT 125.480 264.810 125.860 265.190 ;
      LAYER Metal2 ;
        RECT 125.510 264.750 125.810 271.680 ;
        RECT 126.820 265.350 127.120 271.700 ;
        RECT 128.135 265.380 128.430 272.205 ;
    END
  END s3
  PIN s9_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 134.865 153.085 135.245 153.465 ;
        RECT 131.790 152.590 134.415 153.000 ;
        RECT 133.975 150.150 137.050 150.425 ;
        RECT 133.990 146.725 135.300 147.045 ;
        RECT 131.800 146.170 132.180 146.550 ;
      LAYER Metal2 ;
        RECT 131.840 146.080 132.140 153.020 ;
        RECT 134.050 146.655 134.330 153.015 ;
        RECT 134.900 146.655 135.200 153.475 ;
    END
  END s9_not
  PIN s9
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 127.965 153.095 128.345 153.475 ;
        RECT 125.290 152.670 127.030 152.960 ;
        RECT 126.645 148.075 137.050 148.410 ;
        RECT 126.615 146.755 128.395 147.045 ;
        RECT 125.345 146.140 125.725 146.520 ;
      LAYER Metal2 ;
        RECT 125.375 146.080 125.675 153.010 ;
        RECT 126.685 146.680 126.985 153.030 ;
        RECT 128.000 146.710 128.295 153.535 ;
    END
  END s9
  PIN s4_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 134.920 252.000 135.300 252.380 ;
        RECT 131.845 251.505 134.470 251.915 ;
        RECT 134.030 249.065 137.105 249.340 ;
        RECT 134.045 245.640 135.355 245.960 ;
        RECT 131.855 245.085 132.235 245.465 ;
      LAYER Metal2 ;
        RECT 131.895 244.995 132.195 251.935 ;
        RECT 134.105 245.570 134.385 251.930 ;
        RECT 134.955 245.570 135.255 252.390 ;
    END
  END s4_not
  PIN s4
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 128.020 252.010 128.400 252.390 ;
        RECT 125.345 251.585 127.085 251.875 ;
        RECT 126.700 246.990 137.105 247.325 ;
        RECT 126.670 245.670 128.450 245.960 ;
        RECT 125.400 245.055 125.780 245.435 ;
      LAYER Metal2 ;
        RECT 125.430 244.995 125.730 251.925 ;
        RECT 126.740 245.595 127.040 251.945 ;
        RECT 128.055 245.625 128.350 252.450 ;
    END
  END s4
  PIN s10_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 135.020 133.440 135.400 133.820 ;
        RECT 131.945 132.945 134.570 133.355 ;
        RECT 134.130 130.505 137.205 130.780 ;
        RECT 134.145 127.080 135.455 127.400 ;
        RECT 131.955 126.525 132.335 126.905 ;
      LAYER Metal2 ;
        RECT 131.995 126.435 132.295 133.375 ;
        RECT 134.205 127.010 134.485 133.370 ;
        RECT 135.055 127.010 135.355 133.830 ;
    END
  END s10_not
  PIN s10
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 128.120 133.450 128.500 133.830 ;
        RECT 125.445 133.025 127.185 133.315 ;
        RECT 126.800 128.430 137.205 128.765 ;
        RECT 126.770 127.110 128.550 127.400 ;
        RECT 125.500 126.495 125.880 126.875 ;
      LAYER Metal2 ;
        RECT 125.530 126.435 125.830 133.365 ;
        RECT 126.840 127.035 127.140 133.385 ;
        RECT 128.155 127.065 128.450 133.890 ;
    END
  END s10
  PIN s11_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 135.020 113.645 135.400 114.025 ;
        RECT 131.945 113.150 134.570 113.560 ;
        RECT 134.130 110.710 137.205 110.985 ;
        RECT 134.145 107.285 135.455 107.605 ;
        RECT 131.955 106.730 132.335 107.110 ;
      LAYER Metal2 ;
        RECT 131.995 106.640 132.295 113.580 ;
        RECT 134.205 107.215 134.485 113.575 ;
        RECT 135.055 107.215 135.355 114.035 ;
    END
  END s11_not
  PIN s11
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 128.120 113.655 128.500 114.035 ;
        RECT 125.445 113.230 127.185 113.520 ;
        RECT 126.800 108.635 137.205 108.970 ;
        RECT 126.770 107.315 128.550 107.605 ;
        RECT 125.500 106.700 125.880 107.080 ;
      LAYER Metal2 ;
        RECT 125.530 106.640 125.830 113.570 ;
        RECT 126.840 107.240 127.140 113.590 ;
        RECT 128.155 107.270 128.450 114.095 ;
    END
  END s11
  PIN s12_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 134.940 93.890 135.320 94.270 ;
        RECT 131.865 93.395 134.490 93.805 ;
        RECT 134.050 90.955 137.125 91.230 ;
        RECT 134.065 87.530 135.375 87.850 ;
        RECT 131.875 86.975 132.255 87.355 ;
      LAYER Metal2 ;
        RECT 131.915 86.885 132.215 93.825 ;
        RECT 134.125 87.460 134.405 93.820 ;
        RECT 134.975 87.460 135.275 94.280 ;
    END
  END s12_not
  PIN s12
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 128.040 93.900 128.420 94.280 ;
        RECT 125.365 93.475 127.105 93.765 ;
        RECT 126.720 88.880 137.125 89.215 ;
        RECT 126.690 87.560 128.470 87.850 ;
        RECT 125.420 86.945 125.800 87.325 ;
      LAYER Metal2 ;
        RECT 125.450 86.885 125.750 93.815 ;
        RECT 126.760 87.485 127.060 93.835 ;
        RECT 128.075 87.515 128.370 94.340 ;
    END
  END s12
  PIN s13_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 135.045 74.175 135.425 74.555 ;
        RECT 131.970 73.680 134.595 74.090 ;
        RECT 134.155 71.240 137.230 71.515 ;
        RECT 134.170 67.815 135.480 68.135 ;
        RECT 131.980 67.260 132.360 67.640 ;
      LAYER Metal2 ;
        RECT 132.020 67.170 132.320 74.110 ;
        RECT 134.230 67.745 134.510 74.105 ;
        RECT 135.080 67.745 135.380 74.565 ;
    END
  END s13_not
  PIN s13
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 128.145 74.185 128.525 74.565 ;
        RECT 125.470 73.760 127.210 74.050 ;
        RECT 126.825 69.165 137.230 69.500 ;
        RECT 126.795 67.845 128.575 68.135 ;
        RECT 125.525 67.230 125.905 67.610 ;
      LAYER Metal2 ;
        RECT 125.555 67.170 125.855 74.100 ;
        RECT 126.865 67.770 127.165 74.120 ;
        RECT 128.180 67.800 128.475 74.625 ;
    END
  END s13
  PIN s14_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 135.045 54.205 135.425 54.585 ;
        RECT 131.970 53.710 134.595 54.120 ;
        RECT 134.155 51.270 137.230 51.545 ;
        RECT 134.170 47.845 135.480 48.165 ;
        RECT 131.980 47.290 132.360 47.670 ;
      LAYER Metal2 ;
        RECT 132.020 47.200 132.320 54.140 ;
        RECT 134.230 47.775 134.510 54.135 ;
        RECT 135.080 47.775 135.380 54.595 ;
    END
  END s14_not
  PIN s14
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 128.145 54.215 128.525 54.595 ;
        RECT 125.470 53.790 127.210 54.080 ;
        RECT 126.825 49.195 137.230 49.530 ;
        RECT 126.795 47.875 128.575 48.165 ;
        RECT 125.525 47.260 125.905 47.640 ;
      LAYER Metal2 ;
        RECT 125.555 47.200 125.855 54.130 ;
        RECT 126.865 47.800 127.165 54.150 ;
        RECT 128.180 47.830 128.475 54.655 ;
    END
  END s14
  PIN s15_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 135.045 34.540 135.425 34.920 ;
        RECT 131.970 34.045 134.595 34.455 ;
        RECT 134.155 31.605 137.230 31.880 ;
        RECT 134.170 28.180 135.480 28.500 ;
        RECT 131.980 27.625 132.360 28.005 ;
      LAYER Metal2 ;
        RECT 132.020 27.535 132.320 34.475 ;
        RECT 134.230 28.110 134.510 34.470 ;
        RECT 135.080 28.110 135.380 34.930 ;
    END
  END s15_not
  PIN s15
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 128.145 34.550 128.525 34.930 ;
        RECT 125.470 34.125 127.210 34.415 ;
        RECT 126.825 29.530 137.230 29.865 ;
        RECT 126.795 28.210 128.575 28.500 ;
        RECT 125.525 27.595 125.905 27.975 ;
      LAYER Metal2 ;
        RECT 125.555 27.535 125.855 34.465 ;
        RECT 126.865 28.135 127.165 34.485 ;
        RECT 128.180 28.165 128.475 34.990 ;
    END
  END s15
  PIN z
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 86.780 14.855 87.160 15.235 ;
        RECT 85.180 14.340 86.380 14.630 ;
        RECT 77.445 12.170 86.375 12.470 ;
        RECT 85.970 8.565 87.160 8.850 ;
        RECT 85.190 7.900 85.570 8.280 ;
      LAYER Metal2 ;
        RECT 85.230 7.890 85.530 14.700 ;
        RECT 86.020 8.485 86.330 14.675 ;
        RECT 86.815 8.415 87.115 15.245 ;
    END
  END z
  PIN z_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT 80.320 15.020 83.720 15.455 ;
        RECT 92.100 14.405 92.480 14.785 ;
        RECT 77.415 11.635 83.755 11.905 ;
        RECT 83.330 10.375 89.720 10.665 ;
        RECT 80.310 8.460 80.690 8.840 ;
        RECT 89.310 7.735 92.490 8.055 ;
      LAYER Metal2 ;
        RECT 80.355 8.405 80.655 15.445 ;
        RECT 83.380 10.275 83.700 15.435 ;
        RECT 89.390 7.675 89.670 10.710 ;
        RECT 92.140 7.630 92.440 14.785 ;
    END
  END z_not
  PIN c0_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 112.685 330.930 113.065 331.310 ;
        RECT 110.010 330.505 111.750 330.795 ;
        RECT 123.215 329.745 139.135 330.045 ;
        RECT 124.945 327.090 129.075 327.390 ;
        RECT 131.450 327.040 135.950 327.350 ;
        RECT 111.365 325.910 121.845 326.245 ;
        RECT 111.335 324.590 113.115 324.880 ;
        RECT 110.065 323.975 110.445 324.355 ;
      LAYER Metal2 ;
        RECT 110.095 323.915 110.395 330.845 ;
        RECT 111.405 324.515 111.705 330.865 ;
        RECT 112.720 324.545 113.015 331.370 ;
        RECT 121.405 325.880 121.785 326.260 ;
        RECT 123.255 325.760 123.570 330.085 ;
      LAYER Metal3 ;
        RECT 121.360 325.860 123.645 326.285 ;
    END
  END c0_b
  PIN c0_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 119.585 330.920 119.965 331.300 ;
        RECT 116.510 330.415 119.140 330.870 ;
        RECT 123.750 329.000 140.695 329.300 ;
        RECT 118.695 327.985 121.825 328.260 ;
        RECT 126.175 325.325 129.095 325.625 ;
        RECT 132.640 325.310 136.010 325.610 ;
        RECT 118.710 324.560 120.020 324.880 ;
        RECT 116.520 324.005 116.900 324.385 ;
      LAYER Metal2 ;
        RECT 116.560 323.915 116.860 330.855 ;
        RECT 118.770 324.490 119.050 330.850 ;
        RECT 119.620 324.490 119.920 331.310 ;
        RECT 121.405 327.935 121.785 328.315 ;
        RECT 123.865 327.835 124.145 329.365 ;
        RECT 126.210 325.275 126.510 329.335 ;
        RECT 132.700 325.260 132.980 329.350 ;
      LAYER Metal3 ;
        RECT 121.385 327.935 124.230 328.315 ;
    END
  END c0_not_b
  PIN a0_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 102.885 333.305 104.120 333.685 ;
        RECT 100.860 330.905 104.120 331.285 ;
        RECT 108.290 329.745 121.905 330.045 ;
        RECT 109.485 327.090 113.615 327.390 ;
        RECT 115.990 327.040 120.490 327.350 ;
        RECT 102.745 326.045 106.690 326.380 ;
        RECT 100.840 325.405 104.140 325.785 ;
        RECT 102.655 323.405 104.140 323.785 ;
      LAYER Metal2 ;
        RECT 102.970 323.160 103.285 333.845 ;
        RECT 106.295 326.030 106.675 326.410 ;
        RECT 108.360 326.005 108.670 330.125 ;
        RECT 121.430 329.700 121.725 335.070 ;
      LAYER Metal3 ;
        RECT 121.430 334.615 137.450 335.025 ;
        RECT 106.295 326.020 108.775 326.420 ;
    END
  END a0_b
  PIN a0_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 83.360 333.205 84.560 333.585 ;
        RECT 83.360 330.905 86.620 331.285 ;
        RECT 84.025 328.990 106.580 329.330 ;
        RECT 107.690 329.000 122.335 329.300 ;
        RECT 83.340 325.405 86.640 325.785 ;
        RECT 110.715 325.325 113.635 325.625 ;
        RECT 117.180 325.310 120.550 325.610 ;
        RECT 83.340 323.405 84.625 323.785 ;
      LAYER Metal2 ;
        RECT 84.185 322.675 84.500 333.725 ;
        RECT 106.160 328.920 106.580 329.380 ;
        RECT 107.660 328.915 108.080 329.375 ;
        RECT 110.750 325.275 111.050 329.335 ;
        RECT 117.240 325.260 117.520 329.350 ;
        RECT 122.005 328.870 122.310 334.345 ;
      LAYER Metal3 ;
        RECT 121.960 333.835 137.440 334.290 ;
        RECT 106.130 328.970 108.155 329.355 ;
    END
  END a0_not_b
  PIN a1_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 102.685 313.580 103.920 313.960 ;
        RECT 100.660 311.180 103.920 311.560 ;
        RECT 108.090 310.020 121.705 310.320 ;
        RECT 109.285 307.365 113.415 307.665 ;
        RECT 115.790 307.315 120.290 307.625 ;
        RECT 102.545 306.320 106.490 306.655 ;
        RECT 100.640 305.680 103.940 306.060 ;
        RECT 102.455 303.680 103.940 304.060 ;
      LAYER Metal2 ;
        RECT 102.770 303.435 103.085 314.120 ;
        RECT 106.095 306.305 106.475 306.685 ;
        RECT 108.160 306.280 108.470 310.400 ;
        RECT 121.230 309.975 121.525 315.345 ;
      LAYER Metal3 ;
        RECT 121.230 314.890 137.250 315.300 ;
        RECT 106.095 306.295 108.575 306.695 ;
    END
  END a1_b
  PIN a1_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 83.160 313.480 84.360 313.860 ;
        RECT 83.160 311.180 86.420 311.560 ;
        RECT 83.825 309.265 106.380 309.605 ;
        RECT 107.490 309.275 122.135 309.575 ;
        RECT 83.140 305.680 86.440 306.060 ;
        RECT 110.515 305.600 113.435 305.900 ;
        RECT 116.980 305.585 120.350 305.885 ;
        RECT 83.140 303.680 84.425 304.060 ;
      LAYER Metal2 ;
        RECT 83.985 302.950 84.300 314.000 ;
        RECT 105.960 309.195 106.380 309.655 ;
        RECT 107.460 309.190 107.880 309.650 ;
        RECT 110.550 305.550 110.850 309.610 ;
        RECT 117.040 305.535 117.320 309.625 ;
        RECT 121.805 309.145 122.110 314.620 ;
      LAYER Metal3 ;
        RECT 121.760 314.110 137.240 314.565 ;
        RECT 105.930 309.245 107.955 309.630 ;
    END
  END a1_not_b
  PIN a2_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 102.840 293.935 104.075 294.315 ;
        RECT 100.815 291.535 104.075 291.915 ;
        RECT 108.245 290.375 121.860 290.675 ;
        RECT 109.440 287.720 113.570 288.020 ;
        RECT 115.945 287.670 120.445 287.980 ;
        RECT 102.700 286.675 106.645 287.010 ;
        RECT 100.795 286.035 104.095 286.415 ;
        RECT 102.610 284.035 104.095 284.415 ;
      LAYER Metal2 ;
        RECT 102.925 283.790 103.240 294.475 ;
        RECT 106.250 286.660 106.630 287.040 ;
        RECT 108.315 286.635 108.625 290.755 ;
        RECT 121.385 290.330 121.680 295.700 ;
      LAYER Metal3 ;
        RECT 121.385 295.245 137.405 295.655 ;
        RECT 106.250 286.650 108.730 287.050 ;
    END
  END a2_b
  PIN a2_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 83.315 293.835 84.515 294.215 ;
        RECT 83.315 291.535 86.575 291.915 ;
        RECT 83.980 289.620 106.535 289.960 ;
        RECT 107.645 289.630 122.290 289.930 ;
        RECT 83.295 286.035 86.595 286.415 ;
        RECT 110.670 285.955 113.590 286.255 ;
        RECT 117.135 285.940 120.505 286.240 ;
        RECT 83.295 284.035 84.580 284.415 ;
      LAYER Metal2 ;
        RECT 84.140 283.305 84.455 294.355 ;
        RECT 106.115 289.550 106.535 290.010 ;
        RECT 107.615 289.545 108.035 290.005 ;
        RECT 110.705 285.905 111.005 289.965 ;
        RECT 117.195 285.890 117.475 289.980 ;
        RECT 121.960 289.500 122.265 294.975 ;
      LAYER Metal3 ;
        RECT 121.915 294.465 137.395 294.920 ;
        RECT 106.085 289.600 108.110 289.985 ;
    END
  END a2_not_b
  PIN a3_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 102.840 274.140 104.075 274.520 ;
        RECT 100.815 271.740 104.075 272.120 ;
        RECT 108.245 270.580 121.860 270.880 ;
        RECT 109.440 267.925 113.570 268.225 ;
        RECT 115.945 267.875 120.445 268.185 ;
        RECT 102.700 266.880 106.645 267.215 ;
        RECT 100.795 266.240 104.095 266.620 ;
        RECT 102.610 264.240 104.095 264.620 ;
      LAYER Metal2 ;
        RECT 102.925 263.995 103.240 274.680 ;
        RECT 106.250 266.865 106.630 267.245 ;
        RECT 108.315 266.840 108.625 270.960 ;
        RECT 121.385 270.535 121.680 275.905 ;
      LAYER Metal3 ;
        RECT 121.385 275.450 137.405 275.860 ;
        RECT 106.250 266.855 108.730 267.255 ;
    END
  END a3_b
  PIN a3_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 83.315 274.040 84.515 274.420 ;
        RECT 83.315 271.740 86.575 272.120 ;
        RECT 83.980 269.825 106.535 270.165 ;
        RECT 107.645 269.835 122.290 270.135 ;
        RECT 83.295 266.240 86.595 266.620 ;
        RECT 110.670 266.160 113.590 266.460 ;
        RECT 117.135 266.145 120.505 266.445 ;
        RECT 83.295 264.240 84.580 264.620 ;
      LAYER Metal2 ;
        RECT 84.140 263.510 84.455 274.560 ;
        RECT 106.115 269.755 106.535 270.215 ;
        RECT 107.615 269.750 108.035 270.210 ;
        RECT 110.705 266.110 111.005 270.170 ;
        RECT 117.195 266.095 117.475 270.185 ;
        RECT 121.960 269.705 122.265 275.180 ;
      LAYER Metal3 ;
        RECT 121.915 274.670 137.395 275.125 ;
        RECT 106.085 269.805 108.110 270.190 ;
    END
  END a3_not_b
  PIN a4_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 102.760 254.385 103.995 254.765 ;
        RECT 100.735 251.985 103.995 252.365 ;
        RECT 108.165 250.825 121.780 251.125 ;
        RECT 109.360 248.170 113.490 248.470 ;
        RECT 115.865 248.120 120.365 248.430 ;
        RECT 102.620 247.125 106.565 247.460 ;
        RECT 100.715 246.485 104.015 246.865 ;
        RECT 102.530 244.485 104.015 244.865 ;
      LAYER Metal2 ;
        RECT 102.845 244.240 103.160 254.925 ;
        RECT 106.170 247.110 106.550 247.490 ;
        RECT 108.235 247.085 108.545 251.205 ;
        RECT 121.305 250.780 121.600 256.150 ;
      LAYER Metal3 ;
        RECT 121.305 255.695 137.325 256.105 ;
        RECT 106.170 247.100 108.650 247.500 ;
    END
  END a4_b
  PIN a4_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 83.235 254.285 84.435 254.665 ;
        RECT 83.235 251.985 86.495 252.365 ;
        RECT 83.900 250.070 106.455 250.410 ;
        RECT 107.565 250.080 122.210 250.380 ;
        RECT 83.215 246.485 86.515 246.865 ;
        RECT 110.590 246.405 113.510 246.705 ;
        RECT 117.055 246.390 120.425 246.690 ;
        RECT 83.215 244.485 84.500 244.865 ;
      LAYER Metal2 ;
        RECT 84.060 243.755 84.375 254.805 ;
        RECT 106.035 250.000 106.455 250.460 ;
        RECT 107.535 249.995 107.955 250.455 ;
        RECT 110.625 246.355 110.925 250.415 ;
        RECT 117.115 246.340 117.395 250.430 ;
        RECT 121.880 249.950 122.185 255.425 ;
      LAYER Metal3 ;
        RECT 121.835 254.915 137.315 255.370 ;
        RECT 106.005 250.050 108.030 250.435 ;
    END
  END a4_not_b
  PIN a5_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 102.865 234.670 104.100 235.050 ;
        RECT 100.840 232.270 104.100 232.650 ;
        RECT 108.270 231.110 121.885 231.410 ;
        RECT 109.465 228.455 113.595 228.755 ;
        RECT 115.970 228.405 120.470 228.715 ;
        RECT 102.725 227.410 106.670 227.745 ;
        RECT 100.820 226.770 104.120 227.150 ;
        RECT 102.635 224.770 104.120 225.150 ;
      LAYER Metal2 ;
        RECT 102.950 224.525 103.265 235.210 ;
        RECT 106.275 227.395 106.655 227.775 ;
        RECT 108.340 227.370 108.650 231.490 ;
        RECT 121.410 231.065 121.705 236.435 ;
      LAYER Metal3 ;
        RECT 121.410 235.980 137.430 236.390 ;
        RECT 106.275 227.385 108.755 227.785 ;
    END
  END a5_b
  PIN a5_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 83.340 234.570 84.540 234.950 ;
        RECT 83.340 232.270 86.600 232.650 ;
        RECT 84.005 230.355 106.560 230.695 ;
        RECT 107.670 230.365 122.315 230.665 ;
        RECT 83.320 226.770 86.620 227.150 ;
        RECT 110.695 226.690 113.615 226.990 ;
        RECT 117.160 226.675 120.530 226.975 ;
        RECT 83.320 224.770 84.605 225.150 ;
      LAYER Metal2 ;
        RECT 84.165 224.040 84.480 235.090 ;
        RECT 106.140 230.285 106.560 230.745 ;
        RECT 107.640 230.280 108.060 230.740 ;
        RECT 110.730 226.640 111.030 230.700 ;
        RECT 117.220 226.625 117.500 230.715 ;
        RECT 121.985 230.235 122.290 235.710 ;
      LAYER Metal3 ;
        RECT 121.940 235.200 137.420 235.655 ;
        RECT 106.110 230.335 108.135 230.720 ;
    END
  END a5_not_b
  PIN a6_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 102.865 214.700 104.100 215.080 ;
        RECT 100.840 212.300 104.100 212.680 ;
        RECT 108.270 211.140 121.885 211.440 ;
        RECT 109.465 208.485 113.595 208.785 ;
        RECT 115.970 208.435 120.470 208.745 ;
        RECT 102.725 207.440 106.670 207.775 ;
        RECT 100.820 206.800 104.120 207.180 ;
        RECT 102.635 204.800 104.120 205.180 ;
      LAYER Metal2 ;
        RECT 102.950 204.555 103.265 215.240 ;
        RECT 106.275 207.425 106.655 207.805 ;
        RECT 108.340 207.400 108.650 211.520 ;
        RECT 121.410 211.095 121.705 216.465 ;
      LAYER Metal3 ;
        RECT 121.410 216.010 137.430 216.420 ;
        RECT 106.275 207.415 108.755 207.815 ;
    END
  END a6_b
  PIN a6_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 83.340 214.600 84.540 214.980 ;
        RECT 83.340 212.300 86.600 212.680 ;
        RECT 84.005 210.385 106.560 210.725 ;
        RECT 107.670 210.395 122.315 210.695 ;
        RECT 83.320 206.800 86.620 207.180 ;
        RECT 110.695 206.720 113.615 207.020 ;
        RECT 117.160 206.705 120.530 207.005 ;
        RECT 83.320 204.800 84.605 205.180 ;
      LAYER Metal2 ;
        RECT 84.165 204.070 84.480 215.120 ;
        RECT 106.140 210.315 106.560 210.775 ;
        RECT 107.640 210.310 108.060 210.770 ;
        RECT 110.730 206.670 111.030 210.730 ;
        RECT 117.220 206.655 117.500 210.745 ;
        RECT 121.985 210.265 122.290 215.740 ;
      LAYER Metal3 ;
        RECT 121.940 215.230 137.420 215.685 ;
        RECT 106.110 210.365 108.135 210.750 ;
    END
  END a6_not_b
  PIN a7_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 102.865 195.035 104.100 195.415 ;
        RECT 100.840 192.635 104.100 193.015 ;
        RECT 108.270 191.475 121.885 191.775 ;
        RECT 109.465 188.820 113.595 189.120 ;
        RECT 115.970 188.770 120.470 189.080 ;
        RECT 102.725 187.775 106.670 188.110 ;
        RECT 100.820 187.135 104.120 187.515 ;
        RECT 102.635 185.135 104.120 185.515 ;
      LAYER Metal2 ;
        RECT 102.950 184.890 103.265 195.575 ;
        RECT 106.275 187.760 106.655 188.140 ;
        RECT 108.340 187.735 108.650 191.855 ;
        RECT 121.410 191.430 121.705 196.800 ;
      LAYER Metal3 ;
        RECT 121.410 196.345 137.430 196.755 ;
        RECT 106.275 187.750 108.755 188.150 ;
    END
  END a7_b
  PIN a7_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 83.340 194.935 84.540 195.315 ;
        RECT 83.340 192.635 86.600 193.015 ;
        RECT 84.005 190.720 106.560 191.060 ;
        RECT 107.670 190.730 122.315 191.030 ;
        RECT 83.320 187.135 86.620 187.515 ;
        RECT 110.695 187.055 113.615 187.355 ;
        RECT 117.160 187.040 120.530 187.340 ;
        RECT 83.320 185.135 84.605 185.515 ;
      LAYER Metal2 ;
        RECT 84.165 184.405 84.480 195.455 ;
        RECT 106.140 190.650 106.560 191.110 ;
        RECT 107.640 190.645 108.060 191.105 ;
        RECT 110.730 187.005 111.030 191.065 ;
        RECT 117.220 186.990 117.500 191.080 ;
        RECT 121.985 190.600 122.290 196.075 ;
      LAYER Metal3 ;
        RECT 121.940 195.565 137.420 196.020 ;
        RECT 106.110 190.700 108.135 191.085 ;
    END
  END a7_not_b
  PIN a3_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 42.525 274.020 43.980 274.400 ;
        RECT 42.685 271.720 43.980 272.100 ;
        RECT 56.170 271.720 57.480 272.100 ;
        RECT 41.015 270.395 57.025 270.770 ;
        RECT 10.055 269.815 23.615 270.115 ;
        RECT 25.520 269.815 43.940 270.115 ;
        RECT 12.520 266.140 15.440 266.440 ;
        RECT 18.985 266.125 22.355 266.425 ;
        RECT 27.980 266.140 30.900 266.440 ;
        RECT 34.445 266.125 37.815 266.425 ;
        RECT 42.695 266.220 44.000 266.600 ;
        RECT 56.035 266.220 57.500 266.600 ;
        RECT 42.510 264.220 44.000 264.600 ;
      LAYER Metal2 ;
        RECT 10.055 269.765 10.435 270.145 ;
        RECT 12.555 266.090 12.855 270.150 ;
        RECT 19.045 266.075 19.325 270.165 ;
        RECT 23.235 269.765 23.615 270.145 ;
        RECT 25.505 269.765 25.885 270.170 ;
        RECT 28.015 266.090 28.315 270.150 ;
        RECT 34.505 266.075 34.785 270.165 ;
        RECT 42.815 264.165 43.170 274.470 ;
        RECT 43.480 269.770 43.825 270.825 ;
        RECT 56.325 265.940 56.655 272.135 ;
      LAYER Metal3 ;
        RECT 7.615 269.820 10.460 270.115 ;
        RECT 23.180 269.795 25.920 270.125 ;
    END
  END a3_not_f
  PIN b3
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 17.205 271.785 17.585 272.165 ;
        RECT 15.605 271.270 16.805 271.560 ;
        RECT 10.075 269.100 16.800 269.400 ;
        RECT 16.395 265.495 17.585 265.780 ;
        RECT 15.615 264.830 15.995 265.210 ;
      LAYER Metal2 ;
        RECT 10.100 269.080 10.480 269.460 ;
        RECT 15.655 264.820 15.955 271.630 ;
        RECT 16.445 265.415 16.755 271.605 ;
        RECT 17.240 265.345 17.540 272.175 ;
      LAYER Metal3 ;
        RECT 7.620 269.105 10.495 269.400 ;
    END
  END b3
  PIN b3_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT 10.745 271.985 14.120 272.385 ;
        RECT 22.525 271.335 22.905 271.715 ;
        RECT 10.055 268.480 14.180 268.750 ;
        RECT 13.755 267.305 20.145 267.595 ;
        RECT 10.735 265.390 11.115 265.770 ;
        RECT 19.735 264.665 22.915 264.985 ;
      LAYER Metal2 ;
        RECT 10.065 268.410 10.445 268.790 ;
        RECT 10.780 265.335 11.080 272.375 ;
        RECT 13.805 267.205 14.125 272.365 ;
        RECT 19.815 264.605 20.095 267.640 ;
        RECT 22.565 264.560 22.865 271.715 ;
      LAYER Metal3 ;
        RECT 7.655 268.475 10.450 268.770 ;
    END
  END b3_not
  PIN a4_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 66.090 254.410 67.370 254.790 ;
        RECT 52.590 252.010 53.775 252.390 ;
        RECT 66.090 252.010 67.105 252.390 ;
        RECT 9.930 250.850 23.495 251.165 ;
        RECT 25.385 250.850 39.210 251.150 ;
        RECT 40.885 249.330 67.115 249.720 ;
        RECT 11.160 248.195 15.290 248.495 ;
        RECT 17.665 248.145 22.165 248.455 ;
        RECT 26.620 248.195 30.750 248.495 ;
        RECT 33.125 248.145 37.625 248.455 ;
        RECT 52.570 246.510 53.930 246.890 ;
        RECT 66.070 246.510 67.250 246.890 ;
        RECT 66.070 244.510 67.145 244.890 ;
      LAYER Metal2 ;
        RECT 9.935 250.805 10.315 251.185 ;
        RECT 23.100 250.805 23.480 251.185 ;
        RECT 25.370 250.805 25.750 251.210 ;
        RECT 38.835 250.805 39.195 252.635 ;
        RECT 41.015 249.285 41.430 252.635 ;
        RECT 53.210 252.375 53.520 252.405 ;
        RECT 53.210 246.275 53.525 252.375 ;
        RECT 66.710 244.280 67.040 254.975 ;
      LAYER Metal3 ;
        RECT 38.780 252.250 41.485 252.590 ;
        RECT 7.525 250.845 10.350 251.150 ;
        RECT 23.045 250.835 25.790 251.165 ;
    END
  END a4_f
  PIN a4_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 42.395 254.310 43.850 254.690 ;
        RECT 42.555 252.010 43.850 252.390 ;
        RECT 56.040 252.010 57.350 252.390 ;
        RECT 40.885 250.685 56.895 251.060 ;
        RECT 9.925 250.105 23.485 250.405 ;
        RECT 25.390 250.105 43.810 250.405 ;
        RECT 12.390 246.430 15.310 246.730 ;
        RECT 18.855 246.415 22.225 246.715 ;
        RECT 27.850 246.430 30.770 246.730 ;
        RECT 34.315 246.415 37.685 246.715 ;
        RECT 42.565 246.510 43.870 246.890 ;
        RECT 55.905 246.510 57.370 246.890 ;
        RECT 42.380 244.510 43.870 244.890 ;
      LAYER Metal2 ;
        RECT 9.925 250.055 10.305 250.435 ;
        RECT 12.425 246.380 12.725 250.440 ;
        RECT 18.915 246.365 19.195 250.455 ;
        RECT 23.105 250.055 23.485 250.435 ;
        RECT 25.375 250.055 25.755 250.460 ;
        RECT 27.885 246.380 28.185 250.440 ;
        RECT 34.375 246.365 34.655 250.455 ;
        RECT 42.685 244.455 43.040 254.760 ;
        RECT 43.350 250.060 43.695 251.115 ;
        RECT 56.195 246.230 56.525 252.425 ;
      LAYER Metal3 ;
        RECT 7.485 250.110 10.330 250.405 ;
        RECT 23.050 250.085 25.790 250.415 ;
    END
  END a4_not_f
  PIN b4
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 17.075 252.075 17.455 252.455 ;
        RECT 15.475 251.560 16.675 251.850 ;
        RECT 9.945 249.390 16.670 249.690 ;
        RECT 16.265 245.785 17.455 246.070 ;
        RECT 15.485 245.120 15.865 245.500 ;
      LAYER Metal2 ;
        RECT 9.970 249.370 10.350 249.750 ;
        RECT 15.525 245.110 15.825 251.920 ;
        RECT 16.315 245.705 16.625 251.895 ;
        RECT 17.110 245.635 17.410 252.465 ;
      LAYER Metal3 ;
        RECT 7.490 249.395 10.365 249.690 ;
    END
  END b4
  PIN b4_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT 10.615 252.275 13.990 252.675 ;
        RECT 22.395 251.625 22.775 252.005 ;
        RECT 9.925 248.770 14.050 249.040 ;
        RECT 13.625 247.595 20.015 247.885 ;
        RECT 10.605 245.680 10.985 246.060 ;
        RECT 19.605 244.955 22.785 245.275 ;
      LAYER Metal2 ;
        RECT 9.935 248.700 10.315 249.080 ;
        RECT 10.650 245.625 10.950 252.665 ;
        RECT 13.675 247.495 13.995 252.655 ;
        RECT 19.685 244.895 19.965 247.930 ;
        RECT 22.435 244.850 22.735 252.005 ;
      LAYER Metal3 ;
        RECT 7.525 248.765 10.320 249.060 ;
    END
  END b4_not
  PIN a5_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 66.220 234.650 67.500 235.030 ;
        RECT 52.720 232.250 53.905 232.630 ;
        RECT 66.220 232.250 67.235 232.630 ;
        RECT 10.060 231.090 23.625 231.405 ;
        RECT 25.515 231.090 39.340 231.390 ;
        RECT 41.015 229.570 67.245 229.960 ;
        RECT 11.290 228.435 15.420 228.735 ;
        RECT 17.795 228.385 22.295 228.695 ;
        RECT 26.750 228.435 30.880 228.735 ;
        RECT 33.255 228.385 37.755 228.695 ;
        RECT 52.700 226.750 54.060 227.130 ;
        RECT 66.200 226.750 67.380 227.130 ;
        RECT 66.200 224.750 67.275 225.130 ;
      LAYER Metal2 ;
        RECT 10.065 231.045 10.445 231.425 ;
        RECT 23.230 231.045 23.610 231.425 ;
        RECT 25.500 231.045 25.880 231.450 ;
        RECT 38.965 231.045 39.325 232.875 ;
        RECT 41.145 229.525 41.560 232.875 ;
        RECT 53.340 232.615 53.650 232.645 ;
        RECT 53.340 226.515 53.655 232.615 ;
        RECT 66.840 224.520 67.170 235.215 ;
      LAYER Metal3 ;
        RECT 38.910 232.490 41.615 232.830 ;
        RECT 7.655 231.085 10.480 231.390 ;
        RECT 23.175 231.075 25.920 231.405 ;
    END
  END a5_f
  PIN a5_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 42.525 234.550 43.980 234.930 ;
        RECT 42.685 232.250 43.980 232.630 ;
        RECT 56.170 232.250 57.480 232.630 ;
        RECT 41.015 230.925 57.025 231.300 ;
        RECT 10.055 230.345 23.615 230.645 ;
        RECT 25.520 230.345 43.940 230.645 ;
        RECT 12.520 226.670 15.440 226.970 ;
        RECT 18.985 226.655 22.355 226.955 ;
        RECT 27.980 226.670 30.900 226.970 ;
        RECT 34.445 226.655 37.815 226.955 ;
        RECT 42.695 226.750 44.000 227.130 ;
        RECT 56.035 226.750 57.500 227.130 ;
        RECT 42.510 224.750 44.000 225.130 ;
      LAYER Metal2 ;
        RECT 10.055 230.295 10.435 230.675 ;
        RECT 12.555 226.620 12.855 230.680 ;
        RECT 19.045 226.605 19.325 230.695 ;
        RECT 23.235 230.295 23.615 230.675 ;
        RECT 25.505 230.295 25.885 230.700 ;
        RECT 28.015 226.620 28.315 230.680 ;
        RECT 34.505 226.605 34.785 230.695 ;
        RECT 42.815 224.695 43.170 235.000 ;
        RECT 43.480 230.300 43.825 231.355 ;
        RECT 56.325 226.470 56.655 232.665 ;
      LAYER Metal3 ;
        RECT 7.615 230.350 10.460 230.645 ;
        RECT 23.180 230.325 25.920 230.655 ;
    END
  END a5_not_f
  PIN b5
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 17.205 232.315 17.585 232.695 ;
        RECT 15.605 231.800 16.805 232.090 ;
        RECT 10.075 229.630 16.800 229.930 ;
        RECT 16.395 226.025 17.585 226.310 ;
        RECT 15.615 225.360 15.995 225.740 ;
      LAYER Metal2 ;
        RECT 10.100 229.610 10.480 229.990 ;
        RECT 15.655 225.350 15.955 232.160 ;
        RECT 16.445 225.945 16.755 232.135 ;
        RECT 17.240 225.875 17.540 232.705 ;
      LAYER Metal3 ;
        RECT 7.620 229.635 10.495 229.930 ;
    END
  END b5
  PIN b5_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT 10.745 232.515 14.120 232.915 ;
        RECT 22.525 231.865 22.905 232.245 ;
        RECT 10.055 229.010 14.180 229.280 ;
        RECT 13.755 227.835 20.145 228.125 ;
        RECT 10.735 225.920 11.115 226.300 ;
        RECT 19.735 225.195 22.915 225.515 ;
      LAYER Metal2 ;
        RECT 10.065 228.940 10.445 229.320 ;
        RECT 10.780 225.865 11.080 232.905 ;
        RECT 13.805 227.735 14.125 232.895 ;
        RECT 19.815 225.135 20.095 228.170 ;
        RECT 22.565 225.090 22.865 232.245 ;
      LAYER Metal3 ;
        RECT 7.655 229.005 10.450 229.300 ;
    END
  END b5_not
  PIN a6_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 66.170 214.840 67.450 215.220 ;
        RECT 52.670 212.440 53.855 212.820 ;
        RECT 66.170 212.440 67.185 212.820 ;
        RECT 10.010 211.280 23.575 211.595 ;
        RECT 25.465 211.280 39.290 211.580 ;
        RECT 40.965 209.760 67.195 210.150 ;
        RECT 11.240 208.625 15.370 208.925 ;
        RECT 17.745 208.575 22.245 208.885 ;
        RECT 26.700 208.625 30.830 208.925 ;
        RECT 33.205 208.575 37.705 208.885 ;
        RECT 52.650 206.940 54.010 207.320 ;
        RECT 66.150 206.940 67.330 207.320 ;
        RECT 66.150 204.940 67.225 205.320 ;
      LAYER Metal2 ;
        RECT 10.015 211.235 10.395 211.615 ;
        RECT 23.180 211.235 23.560 211.615 ;
        RECT 25.450 211.235 25.830 211.640 ;
        RECT 38.915 211.235 39.275 213.065 ;
        RECT 41.095 209.715 41.510 213.065 ;
        RECT 53.290 212.805 53.600 212.835 ;
        RECT 53.290 206.705 53.605 212.805 ;
        RECT 66.790 204.710 67.120 215.405 ;
      LAYER Metal3 ;
        RECT 38.860 212.680 41.565 213.020 ;
        RECT 7.605 211.275 10.430 211.580 ;
        RECT 23.125 211.265 25.870 211.595 ;
    END
  END a6_f
  PIN a6_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 42.475 214.740 43.930 215.120 ;
        RECT 42.635 212.440 43.930 212.820 ;
        RECT 56.120 212.440 57.430 212.820 ;
        RECT 40.965 211.115 56.975 211.490 ;
        RECT 10.005 210.535 23.565 210.835 ;
        RECT 25.470 210.535 43.890 210.835 ;
        RECT 12.470 206.860 15.390 207.160 ;
        RECT 18.935 206.845 22.305 207.145 ;
        RECT 27.930 206.860 30.850 207.160 ;
        RECT 34.395 206.845 37.765 207.145 ;
        RECT 42.645 206.940 43.950 207.320 ;
        RECT 55.985 206.940 57.450 207.320 ;
        RECT 42.460 204.940 43.950 205.320 ;
      LAYER Metal2 ;
        RECT 10.005 210.485 10.385 210.865 ;
        RECT 12.505 206.810 12.805 210.870 ;
        RECT 18.995 206.795 19.275 210.885 ;
        RECT 23.185 210.485 23.565 210.865 ;
        RECT 25.455 210.485 25.835 210.890 ;
        RECT 27.965 206.810 28.265 210.870 ;
        RECT 34.455 206.795 34.735 210.885 ;
        RECT 42.765 204.885 43.120 215.190 ;
        RECT 43.430 210.490 43.775 211.545 ;
        RECT 56.275 206.660 56.605 212.855 ;
      LAYER Metal3 ;
        RECT 7.565 210.540 10.410 210.835 ;
        RECT 23.130 210.515 25.870 210.845 ;
    END
  END a6_not_f
  PIN b6
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 17.155 212.505 17.535 212.885 ;
        RECT 15.555 211.990 16.755 212.280 ;
        RECT 10.025 209.820 16.750 210.120 ;
        RECT 16.345 206.215 17.535 206.500 ;
        RECT 15.565 205.550 15.945 205.930 ;
      LAYER Metal2 ;
        RECT 10.050 209.800 10.430 210.180 ;
        RECT 15.605 205.540 15.905 212.350 ;
        RECT 16.395 206.135 16.705 212.325 ;
        RECT 17.190 206.065 17.490 212.895 ;
      LAYER Metal3 ;
        RECT 7.570 209.825 10.445 210.120 ;
    END
  END b6
  PIN b6_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT 10.695 212.705 14.070 213.105 ;
        RECT 22.475 212.055 22.855 212.435 ;
        RECT 10.005 209.200 14.130 209.470 ;
        RECT 13.705 208.025 20.095 208.315 ;
        RECT 10.685 206.110 11.065 206.490 ;
        RECT 19.685 205.385 22.865 205.705 ;
      LAYER Metal2 ;
        RECT 10.015 209.130 10.395 209.510 ;
        RECT 10.730 206.055 11.030 213.095 ;
        RECT 13.755 207.925 14.075 213.085 ;
        RECT 19.765 205.325 20.045 208.360 ;
        RECT 22.515 205.280 22.815 212.435 ;
      LAYER Metal3 ;
        RECT 7.605 209.195 10.400 209.490 ;
    END
  END b6_not
  PIN a7_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 66.140 195.045 67.420 195.425 ;
        RECT 52.640 192.645 53.825 193.025 ;
        RECT 66.140 192.645 67.155 193.025 ;
        RECT 9.980 191.485 23.545 191.800 ;
        RECT 25.435 191.485 39.260 191.785 ;
        RECT 40.935 189.965 67.165 190.355 ;
        RECT 11.210 188.830 15.340 189.130 ;
        RECT 17.715 188.780 22.215 189.090 ;
        RECT 26.670 188.830 30.800 189.130 ;
        RECT 33.175 188.780 37.675 189.090 ;
        RECT 52.620 187.145 53.980 187.525 ;
        RECT 66.120 187.145 67.300 187.525 ;
        RECT 66.120 185.145 67.195 185.525 ;
      LAYER Metal2 ;
        RECT 9.985 191.440 10.365 191.820 ;
        RECT 23.150 191.440 23.530 191.820 ;
        RECT 25.420 191.440 25.800 191.845 ;
        RECT 38.885 191.440 39.245 193.270 ;
        RECT 41.065 189.920 41.480 193.270 ;
        RECT 53.260 193.010 53.570 193.040 ;
        RECT 53.260 186.910 53.575 193.010 ;
        RECT 66.760 184.915 67.090 195.610 ;
      LAYER Metal3 ;
        RECT 38.830 192.885 41.535 193.225 ;
        RECT 7.575 191.480 10.400 191.785 ;
        RECT 23.095 191.470 25.840 191.800 ;
    END
  END a7_f
  PIN a7_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 42.445 194.945 43.900 195.325 ;
        RECT 42.605 192.645 43.900 193.025 ;
        RECT 56.090 192.645 57.400 193.025 ;
        RECT 40.935 191.320 56.945 191.695 ;
        RECT 9.975 190.740 23.535 191.040 ;
        RECT 25.440 190.740 43.860 191.040 ;
        RECT 12.440 187.065 15.360 187.365 ;
        RECT 18.905 187.050 22.275 187.350 ;
        RECT 27.900 187.065 30.820 187.365 ;
        RECT 34.365 187.050 37.735 187.350 ;
        RECT 42.615 187.145 43.920 187.525 ;
        RECT 55.955 187.145 57.420 187.525 ;
        RECT 42.430 185.145 43.920 185.525 ;
      LAYER Metal2 ;
        RECT 9.975 190.690 10.355 191.070 ;
        RECT 12.475 187.015 12.775 191.075 ;
        RECT 18.965 187.000 19.245 191.090 ;
        RECT 23.155 190.690 23.535 191.070 ;
        RECT 25.425 190.690 25.805 191.095 ;
        RECT 27.935 187.015 28.235 191.075 ;
        RECT 34.425 187.000 34.705 191.090 ;
        RECT 42.735 185.090 43.090 195.395 ;
        RECT 43.400 190.695 43.745 191.750 ;
        RECT 56.245 186.865 56.575 193.060 ;
      LAYER Metal3 ;
        RECT 7.535 190.745 10.380 191.040 ;
        RECT 23.100 190.720 25.840 191.050 ;
    END
  END a7_not_f
  PIN b7
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 17.125 192.710 17.505 193.090 ;
        RECT 15.525 192.195 16.725 192.485 ;
        RECT 9.995 190.025 16.720 190.325 ;
        RECT 16.315 186.420 17.505 186.705 ;
        RECT 15.535 185.755 15.915 186.135 ;
      LAYER Metal2 ;
        RECT 10.020 190.005 10.400 190.385 ;
        RECT 15.575 185.745 15.875 192.555 ;
        RECT 16.365 186.340 16.675 192.530 ;
        RECT 17.160 186.270 17.460 193.100 ;
      LAYER Metal3 ;
        RECT 7.540 190.030 10.415 190.325 ;
    END
  END b7
  PIN b7_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT 10.665 192.910 14.040 193.310 ;
        RECT 22.445 192.260 22.825 192.640 ;
        RECT 9.975 189.405 14.100 189.675 ;
        RECT 13.675 188.230 20.065 188.520 ;
        RECT 10.655 186.315 11.035 186.695 ;
        RECT 19.655 185.590 22.835 185.910 ;
      LAYER Metal2 ;
        RECT 9.985 189.335 10.365 189.715 ;
        RECT 10.700 186.260 11.000 193.300 ;
        RECT 13.725 188.130 14.045 193.290 ;
        RECT 19.735 185.530 20.015 188.565 ;
        RECT 22.485 185.485 22.785 192.640 ;
      LAYER Metal3 ;
        RECT 7.575 189.400 10.370 189.695 ;
    END
  END b7_not
  PIN a0_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 66.270 333.360 67.550 333.740 ;
        RECT 52.770 330.960 53.955 331.340 ;
        RECT 66.270 330.960 67.285 331.340 ;
        RECT 10.110 329.800 23.675 330.115 ;
        RECT 25.565 329.800 39.390 330.100 ;
        RECT 41.065 328.280 67.295 328.670 ;
        RECT 11.340 327.145 15.470 327.445 ;
        RECT 17.845 327.095 22.345 327.405 ;
        RECT 26.800 327.145 30.930 327.445 ;
        RECT 33.305 327.095 37.805 327.405 ;
        RECT 52.750 325.460 54.110 325.840 ;
        RECT 66.250 325.460 67.430 325.840 ;
        RECT 66.250 323.460 67.325 323.840 ;
      LAYER Metal2 ;
        RECT 10.115 329.755 10.495 330.135 ;
        RECT 23.280 329.755 23.660 330.135 ;
        RECT 25.550 329.755 25.930 330.160 ;
        RECT 39.015 329.755 39.375 331.585 ;
        RECT 41.195 328.235 41.610 331.585 ;
        RECT 53.390 331.325 53.700 331.355 ;
        RECT 53.390 325.225 53.705 331.325 ;
        RECT 66.890 323.230 67.220 333.925 ;
      LAYER Metal3 ;
        RECT 38.960 331.200 41.665 331.540 ;
        RECT 7.705 329.795 10.530 330.100 ;
        RECT 23.225 329.785 25.970 330.115 ;
    END
  END a0_f
  PIN a0_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 42.575 333.260 44.030 333.640 ;
        RECT 42.735 330.960 44.030 331.340 ;
        RECT 56.220 330.960 57.530 331.340 ;
        RECT 41.065 329.635 57.075 330.010 ;
        RECT 10.105 329.055 23.665 329.355 ;
        RECT 25.570 329.055 43.990 329.355 ;
        RECT 12.570 325.380 15.490 325.680 ;
        RECT 19.035 325.365 22.405 325.665 ;
        RECT 28.030 325.380 30.950 325.680 ;
        RECT 34.495 325.365 37.865 325.665 ;
        RECT 42.745 325.460 44.050 325.840 ;
        RECT 56.085 325.460 57.550 325.840 ;
        RECT 42.560 323.460 44.050 323.840 ;
      LAYER Metal2 ;
        RECT 10.105 329.005 10.485 329.385 ;
        RECT 12.605 325.330 12.905 329.390 ;
        RECT 19.095 325.315 19.375 329.405 ;
        RECT 23.285 329.005 23.665 329.385 ;
        RECT 25.555 329.005 25.935 329.410 ;
        RECT 28.065 325.330 28.365 329.390 ;
        RECT 34.555 325.315 34.835 329.405 ;
        RECT 42.865 323.405 43.220 333.710 ;
        RECT 43.530 329.010 43.875 330.065 ;
        RECT 56.375 325.180 56.705 331.375 ;
      LAYER Metal3 ;
        RECT 7.665 329.060 10.510 329.355 ;
        RECT 23.230 329.035 25.970 329.365 ;
    END
  END a0_not_f
  PIN b0
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 17.255 331.025 17.635 331.405 ;
        RECT 15.655 330.510 16.855 330.800 ;
        RECT 10.125 328.340 16.850 328.640 ;
        RECT 16.445 324.735 17.635 325.020 ;
        RECT 15.665 324.070 16.045 324.450 ;
      LAYER Metal2 ;
        RECT 10.150 328.320 10.530 328.700 ;
        RECT 15.705 324.060 16.005 330.870 ;
        RECT 16.495 324.655 16.805 330.845 ;
        RECT 17.290 324.585 17.590 331.415 ;
      LAYER Metal3 ;
        RECT 7.670 328.345 10.545 328.640 ;
    END
  END b0
  PIN b0_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT 10.795 331.225 14.170 331.625 ;
        RECT 22.575 330.575 22.955 330.955 ;
        RECT 10.105 327.720 14.230 327.990 ;
        RECT 13.805 326.545 20.195 326.835 ;
        RECT 10.785 324.630 11.165 325.010 ;
        RECT 19.785 323.905 22.965 324.225 ;
      LAYER Metal2 ;
        RECT 10.115 327.650 10.495 328.030 ;
        RECT 10.830 324.575 11.130 331.615 ;
        RECT 13.855 326.445 14.175 331.605 ;
        RECT 19.865 323.845 20.145 326.880 ;
        RECT 22.615 323.800 22.915 330.955 ;
      LAYER Metal3 ;
        RECT 7.705 327.715 10.500 328.010 ;
    END
  END b0_not
  PIN a1_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 66.225 313.670 67.505 314.050 ;
        RECT 52.725 311.270 53.910 311.650 ;
        RECT 66.225 311.270 67.240 311.650 ;
        RECT 10.065 310.110 23.630 310.425 ;
        RECT 25.520 310.110 39.345 310.410 ;
        RECT 41.020 308.590 67.250 308.980 ;
        RECT 11.295 307.455 15.425 307.755 ;
        RECT 17.800 307.405 22.300 307.715 ;
        RECT 26.755 307.455 30.885 307.755 ;
        RECT 33.260 307.405 37.760 307.715 ;
        RECT 52.705 305.770 54.065 306.150 ;
        RECT 66.205 305.770 67.385 306.150 ;
        RECT 66.205 303.770 67.280 304.150 ;
      LAYER Metal2 ;
        RECT 10.070 310.065 10.450 310.445 ;
        RECT 23.235 310.065 23.615 310.445 ;
        RECT 25.505 310.065 25.885 310.470 ;
        RECT 38.970 310.065 39.330 311.895 ;
        RECT 41.150 308.545 41.565 311.895 ;
        RECT 53.345 311.635 53.655 311.665 ;
        RECT 53.345 305.535 53.660 311.635 ;
        RECT 66.845 303.540 67.175 314.235 ;
      LAYER Metal3 ;
        RECT 38.915 311.510 41.620 311.850 ;
        RECT 7.660 310.105 10.485 310.410 ;
        RECT 23.180 310.095 25.925 310.425 ;
    END
  END a1_f
  PIN a1_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 42.530 313.570 43.985 313.950 ;
        RECT 42.690 311.270 43.985 311.650 ;
        RECT 56.175 311.270 57.485 311.650 ;
        RECT 41.020 309.945 57.030 310.320 ;
        RECT 10.060 309.365 23.620 309.665 ;
        RECT 25.525 309.365 43.945 309.665 ;
        RECT 12.525 305.690 15.445 305.990 ;
        RECT 18.990 305.675 22.360 305.975 ;
        RECT 27.985 305.690 30.905 305.990 ;
        RECT 34.450 305.675 37.820 305.975 ;
        RECT 42.700 305.770 44.005 306.150 ;
        RECT 56.040 305.770 57.505 306.150 ;
        RECT 42.515 303.770 44.005 304.150 ;
      LAYER Metal2 ;
        RECT 10.060 309.315 10.440 309.695 ;
        RECT 12.560 305.640 12.860 309.700 ;
        RECT 19.050 305.625 19.330 309.715 ;
        RECT 23.240 309.315 23.620 309.695 ;
        RECT 25.510 309.315 25.890 309.720 ;
        RECT 28.020 305.640 28.320 309.700 ;
        RECT 34.510 305.625 34.790 309.715 ;
        RECT 42.820 303.715 43.175 314.020 ;
        RECT 43.485 309.320 43.830 310.375 ;
        RECT 56.330 305.490 56.660 311.685 ;
      LAYER Metal3 ;
        RECT 7.620 309.370 10.465 309.665 ;
        RECT 23.185 309.345 25.925 309.675 ;
    END
  END a1_not_f
  PIN b1
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 17.210 311.335 17.590 311.715 ;
        RECT 15.610 310.820 16.810 311.110 ;
        RECT 10.080 308.650 16.805 308.950 ;
        RECT 16.400 305.045 17.590 305.330 ;
        RECT 15.620 304.380 16.000 304.760 ;
      LAYER Metal2 ;
        RECT 10.105 308.630 10.485 309.010 ;
        RECT 15.660 304.370 15.960 311.180 ;
        RECT 16.450 304.965 16.760 311.155 ;
        RECT 17.245 304.895 17.545 311.725 ;
      LAYER Metal3 ;
        RECT 7.625 308.655 10.500 308.950 ;
    END
  END b1
  PIN b1_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT 10.750 311.535 14.125 311.935 ;
        RECT 22.530 310.885 22.910 311.265 ;
        RECT 10.060 308.030 14.185 308.300 ;
        RECT 13.760 306.855 20.150 307.145 ;
        RECT 10.740 304.940 11.120 305.320 ;
        RECT 19.740 304.215 22.920 304.535 ;
      LAYER Metal2 ;
        RECT 10.070 307.960 10.450 308.340 ;
        RECT 10.785 304.885 11.085 311.925 ;
        RECT 13.810 306.755 14.130 311.915 ;
        RECT 19.820 304.155 20.100 307.190 ;
        RECT 22.570 304.110 22.870 311.265 ;
      LAYER Metal3 ;
        RECT 7.660 308.025 10.455 308.320 ;
    END
  END b1_not
  PIN a2_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 66.415 293.960 67.695 294.340 ;
        RECT 52.915 291.560 54.100 291.940 ;
        RECT 66.415 291.560 67.430 291.940 ;
        RECT 10.255 290.400 23.820 290.715 ;
        RECT 25.710 290.400 39.535 290.700 ;
        RECT 41.210 288.880 67.440 289.270 ;
        RECT 11.485 287.745 15.615 288.045 ;
        RECT 17.990 287.695 22.490 288.005 ;
        RECT 26.945 287.745 31.075 288.045 ;
        RECT 33.450 287.695 37.950 288.005 ;
        RECT 52.895 286.060 54.255 286.440 ;
        RECT 66.395 286.060 67.575 286.440 ;
        RECT 66.395 284.060 67.470 284.440 ;
      LAYER Metal2 ;
        RECT 10.260 290.355 10.640 290.735 ;
        RECT 23.425 290.355 23.805 290.735 ;
        RECT 25.695 290.355 26.075 290.760 ;
        RECT 39.160 290.355 39.520 292.185 ;
        RECT 41.340 288.835 41.755 292.185 ;
        RECT 53.535 291.925 53.845 291.955 ;
        RECT 53.535 285.825 53.850 291.925 ;
        RECT 67.035 283.830 67.365 294.525 ;
      LAYER Metal3 ;
        RECT 39.105 291.800 41.810 292.140 ;
        RECT 7.850 290.395 10.675 290.700 ;
        RECT 23.370 290.385 26.115 290.715 ;
    END
  END a2_f
  PIN a2_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 42.720 293.860 44.175 294.240 ;
        RECT 42.880 291.560 44.175 291.940 ;
        RECT 56.365 291.560 57.675 291.940 ;
        RECT 41.210 290.235 57.220 290.610 ;
        RECT 10.250 289.655 23.810 289.955 ;
        RECT 25.715 289.655 44.135 289.955 ;
        RECT 12.715 285.980 15.635 286.280 ;
        RECT 19.180 285.965 22.550 286.265 ;
        RECT 28.175 285.980 31.095 286.280 ;
        RECT 34.640 285.965 38.010 286.265 ;
        RECT 42.890 286.060 44.195 286.440 ;
        RECT 56.230 286.060 57.695 286.440 ;
        RECT 42.705 284.060 44.195 284.440 ;
      LAYER Metal2 ;
        RECT 10.250 289.605 10.630 289.985 ;
        RECT 12.750 285.930 13.050 289.990 ;
        RECT 19.240 285.915 19.520 290.005 ;
        RECT 23.430 289.605 23.810 289.985 ;
        RECT 25.700 289.605 26.080 290.010 ;
        RECT 28.210 285.930 28.510 289.990 ;
        RECT 34.700 285.915 34.980 290.005 ;
        RECT 43.010 284.005 43.365 294.310 ;
        RECT 43.675 289.610 44.020 290.665 ;
        RECT 56.520 285.780 56.850 291.975 ;
      LAYER Metal3 ;
        RECT 7.810 289.660 10.655 289.955 ;
        RECT 23.375 289.635 26.115 289.965 ;
    END
  END a2_not_f
  PIN b2
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 17.400 291.625 17.780 292.005 ;
        RECT 15.800 291.110 17.000 291.400 ;
        RECT 10.270 288.940 16.995 289.240 ;
        RECT 16.590 285.335 17.780 285.620 ;
        RECT 15.810 284.670 16.190 285.050 ;
      LAYER Metal2 ;
        RECT 10.295 288.920 10.675 289.300 ;
        RECT 15.850 284.660 16.150 291.470 ;
        RECT 16.640 285.255 16.950 291.445 ;
        RECT 17.435 285.185 17.735 292.015 ;
      LAYER Metal3 ;
        RECT 7.815 288.945 10.690 289.240 ;
    END
  END b2
  PIN b2_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT 10.940 291.825 14.315 292.225 ;
        RECT 22.720 291.175 23.100 291.555 ;
        RECT 10.250 288.320 14.375 288.590 ;
        RECT 13.950 287.145 20.340 287.435 ;
        RECT 10.930 285.230 11.310 285.610 ;
        RECT 19.930 284.505 23.110 284.825 ;
      LAYER Metal2 ;
        RECT 10.260 288.250 10.640 288.630 ;
        RECT 10.975 285.175 11.275 292.215 ;
        RECT 14.000 287.045 14.320 292.205 ;
        RECT 20.010 284.445 20.290 287.480 ;
        RECT 22.760 284.400 23.060 291.555 ;
      LAYER Metal3 ;
        RECT 7.850 288.315 10.645 288.610 ;
    END
  END b2_not
  PIN a3_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 66.220 274.120 67.500 274.500 ;
        RECT 52.720 271.720 53.905 272.100 ;
        RECT 66.220 271.720 67.235 272.100 ;
        RECT 10.060 270.560 23.625 270.875 ;
        RECT 25.515 270.560 39.340 270.860 ;
        RECT 41.015 269.040 67.245 269.430 ;
        RECT 11.290 267.905 15.420 268.205 ;
        RECT 17.795 267.855 22.295 268.165 ;
        RECT 26.750 267.905 30.880 268.205 ;
        RECT 33.255 267.855 37.755 268.165 ;
        RECT 52.700 266.220 54.060 266.600 ;
        RECT 66.200 266.220 67.380 266.600 ;
        RECT 66.200 264.220 67.275 264.600 ;
      LAYER Metal2 ;
        RECT 10.065 270.515 10.445 270.895 ;
        RECT 23.230 270.515 23.610 270.895 ;
        RECT 25.500 270.515 25.880 270.920 ;
        RECT 38.965 270.515 39.325 272.345 ;
        RECT 41.145 268.995 41.560 272.345 ;
        RECT 53.340 272.085 53.650 272.115 ;
        RECT 53.340 265.985 53.655 272.085 ;
        RECT 66.840 263.990 67.170 274.685 ;
      LAYER Metal3 ;
        RECT 38.910 271.960 41.615 272.300 ;
        RECT 7.655 270.555 10.480 270.860 ;
        RECT 23.175 270.545 25.920 270.875 ;
    END
  END a3_f
  PIN c0_f
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 32.715 331.025 33.095 331.405 ;
        RECT 31.115 330.510 32.315 330.800 ;
        RECT 25.050 328.340 32.310 328.640 ;
        RECT 31.905 324.735 33.095 325.020 ;
        RECT 31.125 324.070 31.505 324.450 ;
      LAYER Metal2 ;
        RECT 25.070 326.570 25.390 328.700 ;
        RECT 31.165 324.060 31.465 330.870 ;
        RECT 31.955 324.655 32.265 330.845 ;
        RECT 32.750 324.585 33.050 331.415 ;
      LAYER Metal3 ;
        RECT 4.750 326.640 25.455 326.935 ;
    END
  END c0_f
  PIN c0_f_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT 26.255 331.185 29.660 331.625 ;
        RECT 38.035 330.575 38.415 330.955 ;
        RECT 25.605 327.805 29.690 328.075 ;
        RECT 29.265 326.545 35.655 326.835 ;
        RECT 26.245 324.630 26.625 325.010 ;
        RECT 35.245 323.905 38.425 324.225 ;
      LAYER Metal2 ;
        RECT 25.680 325.730 25.960 328.135 ;
        RECT 26.290 324.575 26.590 331.615 ;
        RECT 29.315 326.445 29.640 331.605 ;
        RECT 35.325 323.845 35.605 326.880 ;
        RECT 38.075 323.800 38.375 330.955 ;
      LAYER Metal3 ;
        RECT 4.570 325.775 26.040 326.070 ;
    END
  END c0_f_not
  PIN b12_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT 10.635 94.165 14.010 94.565 ;
        RECT 22.415 93.515 22.795 93.895 ;
        RECT 9.945 90.660 14.070 90.930 ;
        RECT 13.645 89.485 20.035 89.775 ;
        RECT 10.625 87.570 11.005 87.950 ;
        RECT 19.625 86.845 22.805 87.165 ;
      LAYER Metal2 ;
        RECT 9.955 90.590 10.335 90.970 ;
        RECT 10.670 87.515 10.970 94.555 ;
        RECT 13.695 89.385 14.015 94.545 ;
        RECT 19.705 86.785 19.985 89.820 ;
        RECT 22.455 86.740 22.755 93.895 ;
      LAYER Metal3 ;
        RECT 7.545 90.655 10.340 90.950 ;
    END
  END b12_not
  PIN a13_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 66.240 76.540 67.520 76.920 ;
        RECT 52.740 74.140 53.925 74.520 ;
        RECT 66.240 74.140 67.255 74.520 ;
        RECT 10.080 72.980 23.645 73.295 ;
        RECT 25.535 72.980 39.360 73.280 ;
        RECT 41.035 71.460 67.265 71.850 ;
        RECT 11.310 70.325 15.440 70.625 ;
        RECT 17.815 70.275 22.315 70.585 ;
        RECT 26.770 70.325 30.900 70.625 ;
        RECT 33.275 70.275 37.775 70.585 ;
        RECT 52.720 68.640 54.080 69.020 ;
        RECT 66.220 68.640 67.400 69.020 ;
        RECT 66.220 66.640 67.295 67.020 ;
      LAYER Metal2 ;
        RECT 10.085 72.935 10.465 73.315 ;
        RECT 23.250 72.935 23.630 73.315 ;
        RECT 25.520 72.935 25.900 73.340 ;
        RECT 38.985 72.935 39.345 74.765 ;
        RECT 41.165 71.415 41.580 74.765 ;
        RECT 53.360 74.505 53.670 74.535 ;
        RECT 53.360 68.405 53.675 74.505 ;
        RECT 66.860 66.410 67.190 77.105 ;
      LAYER Metal3 ;
        RECT 38.930 74.380 41.635 74.720 ;
        RECT 7.675 72.975 10.500 73.280 ;
        RECT 23.195 72.965 25.940 73.295 ;
    END
  END a13_f
  PIN a13_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 42.545 76.440 44.000 76.820 ;
        RECT 42.705 74.140 44.000 74.520 ;
        RECT 56.190 74.140 57.500 74.520 ;
        RECT 41.035 72.815 57.045 73.190 ;
        RECT 10.075 72.235 23.635 72.535 ;
        RECT 25.540 72.235 43.960 72.535 ;
        RECT 12.540 68.560 15.460 68.860 ;
        RECT 19.005 68.545 22.375 68.845 ;
        RECT 28.000 68.560 30.920 68.860 ;
        RECT 34.465 68.545 37.835 68.845 ;
        RECT 42.715 68.640 44.020 69.020 ;
        RECT 56.055 68.640 57.520 69.020 ;
        RECT 42.530 66.640 44.020 67.020 ;
      LAYER Metal2 ;
        RECT 10.075 72.185 10.455 72.565 ;
        RECT 12.575 68.510 12.875 72.570 ;
        RECT 19.065 68.495 19.345 72.585 ;
        RECT 23.255 72.185 23.635 72.565 ;
        RECT 25.525 72.185 25.905 72.590 ;
        RECT 28.035 68.510 28.335 72.570 ;
        RECT 34.525 68.495 34.805 72.585 ;
        RECT 42.835 66.585 43.190 76.890 ;
        RECT 43.500 72.190 43.845 73.245 ;
        RECT 56.345 68.360 56.675 74.555 ;
      LAYER Metal3 ;
        RECT 7.635 72.240 10.480 72.535 ;
        RECT 23.200 72.215 25.940 72.545 ;
    END
  END a13_not_f
  PIN b13
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 17.225 74.205 17.605 74.585 ;
        RECT 15.625 73.690 16.825 73.980 ;
        RECT 10.095 71.520 16.820 71.820 ;
        RECT 16.415 67.915 17.605 68.200 ;
        RECT 15.635 67.250 16.015 67.630 ;
      LAYER Metal2 ;
        RECT 10.120 71.500 10.500 71.880 ;
        RECT 15.675 67.240 15.975 74.050 ;
        RECT 16.465 67.835 16.775 74.025 ;
        RECT 17.260 67.765 17.560 74.595 ;
      LAYER Metal3 ;
        RECT 7.640 71.525 10.515 71.820 ;
    END
  END b13
  PIN b13_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT 10.765 74.405 14.140 74.805 ;
        RECT 22.545 73.755 22.925 74.135 ;
        RECT 10.075 70.900 14.200 71.170 ;
        RECT 13.775 69.725 20.165 70.015 ;
        RECT 10.755 67.810 11.135 68.190 ;
        RECT 19.755 67.085 22.935 67.405 ;
      LAYER Metal2 ;
        RECT 10.085 70.830 10.465 71.210 ;
        RECT 10.800 67.755 11.100 74.795 ;
        RECT 13.825 69.625 14.145 74.785 ;
        RECT 19.835 67.025 20.115 70.060 ;
        RECT 22.585 66.980 22.885 74.135 ;
      LAYER Metal3 ;
        RECT 7.675 70.895 10.470 71.190 ;
    END
  END b13_not
  PIN a14_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 66.190 56.730 67.470 57.110 ;
        RECT 52.690 54.330 53.875 54.710 ;
        RECT 66.190 54.330 67.205 54.710 ;
        RECT 10.030 53.170 23.595 53.485 ;
        RECT 25.485 53.170 39.310 53.470 ;
        RECT 40.985 51.650 67.215 52.040 ;
        RECT 11.260 50.515 15.390 50.815 ;
        RECT 17.765 50.465 22.265 50.775 ;
        RECT 26.720 50.515 30.850 50.815 ;
        RECT 33.225 50.465 37.725 50.775 ;
        RECT 52.670 48.830 54.030 49.210 ;
        RECT 66.170 48.830 67.350 49.210 ;
        RECT 66.170 46.830 67.245 47.210 ;
      LAYER Metal2 ;
        RECT 10.035 53.125 10.415 53.505 ;
        RECT 23.200 53.125 23.580 53.505 ;
        RECT 25.470 53.125 25.850 53.530 ;
        RECT 38.935 53.125 39.295 54.955 ;
        RECT 41.115 51.605 41.530 54.955 ;
        RECT 53.310 54.695 53.620 54.725 ;
        RECT 53.310 48.595 53.625 54.695 ;
        RECT 66.810 46.600 67.140 57.295 ;
      LAYER Metal3 ;
        RECT 38.880 54.570 41.585 54.910 ;
        RECT 7.625 53.165 10.450 53.470 ;
        RECT 23.145 53.155 25.890 53.485 ;
    END
  END a14_f
  PIN a14_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 42.495 56.630 43.950 57.010 ;
        RECT 42.655 54.330 43.950 54.710 ;
        RECT 56.140 54.330 57.450 54.710 ;
        RECT 40.985 53.005 56.995 53.380 ;
        RECT 10.025 52.425 23.585 52.725 ;
        RECT 25.490 52.425 43.910 52.725 ;
        RECT 12.490 48.750 15.410 49.050 ;
        RECT 18.955 48.735 22.325 49.035 ;
        RECT 27.950 48.750 30.870 49.050 ;
        RECT 34.415 48.735 37.785 49.035 ;
        RECT 42.665 48.830 43.970 49.210 ;
        RECT 56.005 48.830 57.470 49.210 ;
        RECT 42.480 46.830 43.970 47.210 ;
      LAYER Metal2 ;
        RECT 10.025 52.375 10.405 52.755 ;
        RECT 12.525 48.700 12.825 52.760 ;
        RECT 19.015 48.685 19.295 52.775 ;
        RECT 23.205 52.375 23.585 52.755 ;
        RECT 25.475 52.375 25.855 52.780 ;
        RECT 27.985 48.700 28.285 52.760 ;
        RECT 34.475 48.685 34.755 52.775 ;
        RECT 42.785 46.775 43.140 57.080 ;
        RECT 43.450 52.380 43.795 53.435 ;
        RECT 56.295 48.550 56.625 54.745 ;
      LAYER Metal3 ;
        RECT 7.585 52.430 10.430 52.725 ;
        RECT 23.150 52.405 25.890 52.735 ;
    END
  END a14_not_f
  PIN b14
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 17.175 54.395 17.555 54.775 ;
        RECT 15.575 53.880 16.775 54.170 ;
        RECT 10.045 51.710 16.770 52.010 ;
        RECT 16.365 48.105 17.555 48.390 ;
        RECT 15.585 47.440 15.965 47.820 ;
      LAYER Metal2 ;
        RECT 10.070 51.690 10.450 52.070 ;
        RECT 15.625 47.430 15.925 54.240 ;
        RECT 16.415 48.025 16.725 54.215 ;
        RECT 17.210 47.955 17.510 54.785 ;
      LAYER Metal3 ;
        RECT 7.590 51.715 10.465 52.010 ;
    END
  END b14
  PIN b14_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT 10.715 54.595 14.090 54.995 ;
        RECT 22.495 53.945 22.875 54.325 ;
        RECT 10.025 51.090 14.150 51.360 ;
        RECT 13.725 49.915 20.115 50.205 ;
        RECT 10.705 48.000 11.085 48.380 ;
        RECT 19.705 47.275 22.885 47.595 ;
      LAYER Metal2 ;
        RECT 10.035 51.020 10.415 51.400 ;
        RECT 10.750 47.945 11.050 54.985 ;
        RECT 13.775 49.815 14.095 54.975 ;
        RECT 19.785 47.215 20.065 50.250 ;
        RECT 22.535 47.170 22.835 54.325 ;
      LAYER Metal3 ;
        RECT 7.625 51.085 10.420 51.380 ;
    END
  END b14_not
  PIN a15_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 66.160 36.935 67.440 37.315 ;
        RECT 52.660 34.535 53.845 34.915 ;
        RECT 66.160 34.535 67.175 34.915 ;
        RECT 10.000 33.375 23.565 33.690 ;
        RECT 25.455 33.375 39.280 33.675 ;
        RECT 40.955 31.855 67.185 32.245 ;
        RECT 11.230 30.720 15.360 31.020 ;
        RECT 17.735 30.670 22.235 30.980 ;
        RECT 26.690 30.720 30.820 31.020 ;
        RECT 33.195 30.670 37.695 30.980 ;
        RECT 52.640 29.035 54.000 29.415 ;
        RECT 66.140 29.035 67.320 29.415 ;
        RECT 66.140 27.035 67.215 27.415 ;
      LAYER Metal2 ;
        RECT 10.005 33.330 10.385 33.710 ;
        RECT 23.170 33.330 23.550 33.710 ;
        RECT 25.440 33.330 25.820 33.735 ;
        RECT 38.905 33.330 39.265 35.160 ;
        RECT 41.085 31.810 41.500 35.160 ;
        RECT 53.280 34.900 53.590 34.930 ;
        RECT 53.280 28.800 53.595 34.900 ;
        RECT 66.780 26.805 67.110 37.500 ;
      LAYER Metal3 ;
        RECT 38.850 34.775 41.555 35.115 ;
        RECT 7.595 33.370 10.420 33.675 ;
        RECT 23.115 33.360 25.860 33.690 ;
    END
  END a15_f
  PIN a15_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 42.465 36.835 43.920 37.215 ;
        RECT 42.625 34.535 43.920 34.915 ;
        RECT 56.110 34.535 57.420 34.915 ;
        RECT 40.955 33.210 56.965 33.585 ;
        RECT 9.995 32.630 23.555 32.930 ;
        RECT 25.460 32.630 43.880 32.930 ;
        RECT 12.460 28.955 15.380 29.255 ;
        RECT 18.925 28.940 22.295 29.240 ;
        RECT 27.920 28.955 30.840 29.255 ;
        RECT 34.385 28.940 37.755 29.240 ;
        RECT 42.635 29.035 43.940 29.415 ;
        RECT 55.975 29.035 57.440 29.415 ;
        RECT 42.450 27.035 43.940 27.415 ;
      LAYER Metal2 ;
        RECT 9.995 32.580 10.375 32.960 ;
        RECT 12.495 28.905 12.795 32.965 ;
        RECT 18.985 28.890 19.265 32.980 ;
        RECT 23.175 32.580 23.555 32.960 ;
        RECT 25.445 32.580 25.825 32.985 ;
        RECT 27.955 28.905 28.255 32.965 ;
        RECT 34.445 28.890 34.725 32.980 ;
        RECT 42.755 26.980 43.110 37.285 ;
        RECT 43.420 32.585 43.765 33.640 ;
        RECT 56.265 28.755 56.595 34.950 ;
      LAYER Metal3 ;
        RECT 7.555 32.635 10.400 32.930 ;
        RECT 23.120 32.610 25.860 32.940 ;
    END
  END a15_not_f
  PIN b15
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 17.145 34.600 17.525 34.980 ;
        RECT 15.545 34.085 16.745 34.375 ;
        RECT 10.015 31.915 16.740 32.215 ;
        RECT 16.335 28.310 17.525 28.595 ;
        RECT 15.555 27.645 15.935 28.025 ;
      LAYER Metal2 ;
        RECT 10.040 31.895 10.420 32.275 ;
        RECT 15.595 27.635 15.895 34.445 ;
        RECT 16.385 28.230 16.695 34.420 ;
        RECT 17.180 28.160 17.480 34.990 ;
      LAYER Metal3 ;
        RECT 7.560 31.920 10.435 32.215 ;
    END
  END b15
  PIN b15_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT 10.685 34.800 14.060 35.200 ;
        RECT 22.465 34.150 22.845 34.530 ;
        RECT 9.995 31.295 14.120 31.565 ;
        RECT 13.695 30.120 20.085 30.410 ;
        RECT 10.675 28.205 11.055 28.585 ;
        RECT 19.675 27.480 22.855 27.800 ;
      LAYER Metal2 ;
        RECT 10.005 31.225 10.385 31.605 ;
        RECT 10.720 28.150 11.020 35.190 ;
        RECT 13.745 30.020 14.065 35.180 ;
        RECT 19.755 27.420 20.035 30.455 ;
        RECT 22.505 27.375 22.805 34.530 ;
      LAYER Metal3 ;
        RECT 7.595 31.290 10.390 31.585 ;
    END
  END b15_not
  PIN a8_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 66.290 175.250 67.570 175.630 ;
        RECT 52.790 172.850 53.975 173.230 ;
        RECT 66.290 172.850 67.305 173.230 ;
        RECT 10.130 171.690 23.695 172.005 ;
        RECT 25.585 171.690 39.410 171.990 ;
        RECT 41.085 170.170 67.315 170.560 ;
        RECT 11.360 169.035 15.490 169.335 ;
        RECT 17.865 168.985 22.365 169.295 ;
        RECT 26.820 169.035 30.950 169.335 ;
        RECT 33.325 168.985 37.825 169.295 ;
        RECT 52.770 167.350 54.130 167.730 ;
        RECT 66.270 167.350 67.450 167.730 ;
        RECT 66.270 165.350 67.345 165.730 ;
      LAYER Metal2 ;
        RECT 10.135 171.645 10.515 172.025 ;
        RECT 23.300 171.645 23.680 172.025 ;
        RECT 25.570 171.645 25.950 172.050 ;
        RECT 39.035 171.645 39.395 173.475 ;
        RECT 41.215 170.125 41.630 173.475 ;
        RECT 53.410 173.215 53.720 173.245 ;
        RECT 53.410 167.115 53.725 173.215 ;
        RECT 66.910 165.120 67.240 175.815 ;
      LAYER Metal3 ;
        RECT 38.980 173.090 41.685 173.430 ;
        RECT 7.725 171.685 10.550 171.990 ;
        RECT 23.245 171.675 25.990 172.005 ;
    END
  END a8_f
  PIN a8_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 42.595 175.150 44.050 175.530 ;
        RECT 42.755 172.850 44.050 173.230 ;
        RECT 56.240 172.850 57.550 173.230 ;
        RECT 41.085 171.525 57.095 171.900 ;
        RECT 10.125 170.945 23.685 171.245 ;
        RECT 25.590 170.945 44.010 171.245 ;
        RECT 12.590 167.270 15.510 167.570 ;
        RECT 19.055 167.255 22.425 167.555 ;
        RECT 28.050 167.270 30.970 167.570 ;
        RECT 34.515 167.255 37.885 167.555 ;
        RECT 42.765 167.350 44.070 167.730 ;
        RECT 56.105 167.350 57.570 167.730 ;
        RECT 42.580 165.350 44.070 165.730 ;
      LAYER Metal2 ;
        RECT 10.125 170.895 10.505 171.275 ;
        RECT 12.625 167.220 12.925 171.280 ;
        RECT 19.115 167.205 19.395 171.295 ;
        RECT 23.305 170.895 23.685 171.275 ;
        RECT 25.575 170.895 25.955 171.300 ;
        RECT 28.085 167.220 28.385 171.280 ;
        RECT 34.575 167.205 34.855 171.295 ;
        RECT 42.885 165.295 43.240 175.600 ;
        RECT 43.550 170.900 43.895 171.955 ;
        RECT 56.395 167.070 56.725 173.265 ;
      LAYER Metal3 ;
        RECT 7.685 170.950 10.530 171.245 ;
        RECT 23.250 170.925 25.990 171.255 ;
    END
  END a8_not_f
  PIN b8
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 17.275 172.915 17.655 173.295 ;
        RECT 15.675 172.400 16.875 172.690 ;
        RECT 10.145 170.230 16.870 170.530 ;
        RECT 16.465 166.625 17.655 166.910 ;
        RECT 15.685 165.960 16.065 166.340 ;
      LAYER Metal2 ;
        RECT 10.170 170.210 10.550 170.590 ;
        RECT 15.725 165.950 16.025 172.760 ;
        RECT 16.515 166.545 16.825 172.735 ;
        RECT 17.310 166.475 17.610 173.305 ;
      LAYER Metal3 ;
        RECT 7.690 170.235 10.565 170.530 ;
    END
  END b8
  PIN b8_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT 10.815 173.115 14.190 173.515 ;
        RECT 22.595 172.465 22.975 172.845 ;
        RECT 10.125 169.610 14.250 169.880 ;
        RECT 13.825 168.435 20.215 168.725 ;
        RECT 10.805 166.520 11.185 166.900 ;
        RECT 19.805 165.795 22.985 166.115 ;
      LAYER Metal2 ;
        RECT 10.135 169.540 10.515 169.920 ;
        RECT 10.850 166.465 11.150 173.505 ;
        RECT 13.875 168.335 14.195 173.495 ;
        RECT 19.885 165.735 20.165 168.770 ;
        RECT 22.635 165.690 22.935 172.845 ;
      LAYER Metal3 ;
        RECT 7.725 169.605 10.520 169.900 ;
    END
  END b8_not
  PIN a9_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 66.245 155.560 67.525 155.940 ;
        RECT 52.745 153.160 53.930 153.540 ;
        RECT 66.245 153.160 67.260 153.540 ;
        RECT 10.085 152.000 23.650 152.315 ;
        RECT 25.540 152.000 39.365 152.300 ;
        RECT 41.040 150.480 67.270 150.870 ;
        RECT 11.315 149.345 15.445 149.645 ;
        RECT 17.820 149.295 22.320 149.605 ;
        RECT 26.775 149.345 30.905 149.645 ;
        RECT 33.280 149.295 37.780 149.605 ;
        RECT 52.725 147.660 54.085 148.040 ;
        RECT 66.225 147.660 67.405 148.040 ;
        RECT 66.225 145.660 67.300 146.040 ;
      LAYER Metal2 ;
        RECT 10.090 151.955 10.470 152.335 ;
        RECT 23.255 151.955 23.635 152.335 ;
        RECT 25.525 151.955 25.905 152.360 ;
        RECT 38.990 151.955 39.350 153.785 ;
        RECT 41.170 150.435 41.585 153.785 ;
        RECT 53.365 153.525 53.675 153.555 ;
        RECT 53.365 147.425 53.680 153.525 ;
        RECT 66.865 145.430 67.195 156.125 ;
      LAYER Metal3 ;
        RECT 38.935 153.400 41.640 153.740 ;
        RECT 7.680 151.995 10.505 152.300 ;
        RECT 23.200 151.985 25.945 152.315 ;
    END
  END a9_f
  PIN a9_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 42.550 155.460 44.005 155.840 ;
        RECT 42.710 153.160 44.005 153.540 ;
        RECT 56.195 153.160 57.505 153.540 ;
        RECT 41.040 151.835 57.050 152.210 ;
        RECT 10.080 151.255 23.640 151.555 ;
        RECT 25.545 151.255 43.965 151.555 ;
        RECT 12.545 147.580 15.465 147.880 ;
        RECT 19.010 147.565 22.380 147.865 ;
        RECT 28.005 147.580 30.925 147.880 ;
        RECT 34.470 147.565 37.840 147.865 ;
        RECT 42.720 147.660 44.025 148.040 ;
        RECT 56.060 147.660 57.525 148.040 ;
        RECT 42.535 145.660 44.025 146.040 ;
      LAYER Metal2 ;
        RECT 10.080 151.205 10.460 151.585 ;
        RECT 12.580 147.530 12.880 151.590 ;
        RECT 19.070 147.515 19.350 151.605 ;
        RECT 23.260 151.205 23.640 151.585 ;
        RECT 25.530 151.205 25.910 151.610 ;
        RECT 28.040 147.530 28.340 151.590 ;
        RECT 34.530 147.515 34.810 151.605 ;
        RECT 42.840 145.605 43.195 155.910 ;
        RECT 43.505 151.210 43.850 152.265 ;
        RECT 56.350 147.380 56.680 153.575 ;
      LAYER Metal3 ;
        RECT 7.640 151.260 10.485 151.555 ;
        RECT 23.205 151.235 25.945 151.565 ;
    END
  END a9_not_f
  PIN b9
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 17.230 153.225 17.610 153.605 ;
        RECT 15.630 152.710 16.830 153.000 ;
        RECT 10.100 150.540 16.825 150.840 ;
        RECT 16.420 146.935 17.610 147.220 ;
        RECT 15.640 146.270 16.020 146.650 ;
      LAYER Metal2 ;
        RECT 10.125 150.520 10.505 150.900 ;
        RECT 15.680 146.260 15.980 153.070 ;
        RECT 16.470 146.855 16.780 153.045 ;
        RECT 17.265 146.785 17.565 153.615 ;
      LAYER Metal3 ;
        RECT 7.645 150.545 10.520 150.840 ;
    END
  END b9
  PIN b9_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT 10.770 153.425 14.145 153.825 ;
        RECT 22.550 152.775 22.930 153.155 ;
        RECT 10.080 149.920 14.205 150.190 ;
        RECT 13.780 148.745 20.170 149.035 ;
        RECT 10.760 146.830 11.140 147.210 ;
        RECT 19.760 146.105 22.940 146.425 ;
      LAYER Metal2 ;
        RECT 10.090 149.850 10.470 150.230 ;
        RECT 10.805 146.775 11.105 153.815 ;
        RECT 13.830 148.645 14.150 153.805 ;
        RECT 19.840 146.045 20.120 149.080 ;
        RECT 22.590 146.000 22.890 153.155 ;
      LAYER Metal3 ;
        RECT 7.680 149.915 10.475 150.210 ;
    END
  END b9_not
  PIN a10_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 66.435 135.850 67.715 136.230 ;
        RECT 52.935 133.450 54.120 133.830 ;
        RECT 66.435 133.450 67.450 133.830 ;
        RECT 10.275 132.290 23.840 132.605 ;
        RECT 25.730 132.290 39.555 132.590 ;
        RECT 41.230 130.770 67.460 131.160 ;
        RECT 11.505 129.635 15.635 129.935 ;
        RECT 18.010 129.585 22.510 129.895 ;
        RECT 26.965 129.635 31.095 129.935 ;
        RECT 33.470 129.585 37.970 129.895 ;
        RECT 52.915 127.950 54.275 128.330 ;
        RECT 66.415 127.950 67.595 128.330 ;
        RECT 66.415 125.950 67.490 126.330 ;
      LAYER Metal2 ;
        RECT 10.280 132.245 10.660 132.625 ;
        RECT 23.445 132.245 23.825 132.625 ;
        RECT 25.715 132.245 26.095 132.650 ;
        RECT 39.180 132.245 39.540 134.075 ;
        RECT 41.360 130.725 41.775 134.075 ;
        RECT 53.555 133.815 53.865 133.845 ;
        RECT 53.555 127.715 53.870 133.815 ;
        RECT 67.055 125.720 67.385 136.415 ;
      LAYER Metal3 ;
        RECT 39.125 133.690 41.830 134.030 ;
        RECT 7.870 132.285 10.695 132.590 ;
        RECT 23.390 132.275 26.135 132.605 ;
    END
  END a10_f
  PIN a10_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 42.740 135.750 44.195 136.130 ;
        RECT 42.900 133.450 44.195 133.830 ;
        RECT 56.385 133.450 57.695 133.830 ;
        RECT 41.230 132.125 57.240 132.500 ;
        RECT 10.270 131.545 23.830 131.845 ;
        RECT 25.735 131.545 44.155 131.845 ;
        RECT 12.735 127.870 15.655 128.170 ;
        RECT 19.200 127.855 22.570 128.155 ;
        RECT 28.195 127.870 31.115 128.170 ;
        RECT 34.660 127.855 38.030 128.155 ;
        RECT 42.910 127.950 44.215 128.330 ;
        RECT 56.250 127.950 57.715 128.330 ;
        RECT 42.725 125.950 44.215 126.330 ;
      LAYER Metal2 ;
        RECT 10.270 131.495 10.650 131.875 ;
        RECT 12.770 127.820 13.070 131.880 ;
        RECT 19.260 127.805 19.540 131.895 ;
        RECT 23.450 131.495 23.830 131.875 ;
        RECT 25.720 131.495 26.100 131.900 ;
        RECT 28.230 127.820 28.530 131.880 ;
        RECT 34.720 127.805 35.000 131.895 ;
        RECT 43.030 125.895 43.385 136.200 ;
        RECT 43.695 131.500 44.040 132.555 ;
        RECT 56.540 127.670 56.870 133.865 ;
      LAYER Metal3 ;
        RECT 7.830 131.550 10.675 131.845 ;
        RECT 23.395 131.525 26.135 131.855 ;
    END
  END a10_not_f
  PIN b10
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 17.420 133.515 17.800 133.895 ;
        RECT 15.820 133.000 17.020 133.290 ;
        RECT 10.290 130.830 17.015 131.130 ;
        RECT 16.610 127.225 17.800 127.510 ;
        RECT 15.830 126.560 16.210 126.940 ;
      LAYER Metal2 ;
        RECT 10.315 130.810 10.695 131.190 ;
        RECT 15.870 126.550 16.170 133.360 ;
        RECT 16.660 127.145 16.970 133.335 ;
        RECT 17.455 127.075 17.755 133.905 ;
      LAYER Metal3 ;
        RECT 7.835 130.835 10.710 131.130 ;
    END
  END b10
  PIN b10_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT 10.960 133.715 14.335 134.115 ;
        RECT 22.740 133.065 23.120 133.445 ;
        RECT 10.270 130.210 14.395 130.480 ;
        RECT 13.970 129.035 20.360 129.325 ;
        RECT 10.950 127.120 11.330 127.500 ;
        RECT 19.950 126.395 23.130 126.715 ;
      LAYER Metal2 ;
        RECT 10.280 130.140 10.660 130.520 ;
        RECT 10.995 127.065 11.295 134.105 ;
        RECT 14.020 128.935 14.340 134.095 ;
        RECT 20.030 126.335 20.310 129.370 ;
        RECT 22.780 126.290 23.080 133.445 ;
      LAYER Metal3 ;
        RECT 7.870 130.205 10.665 130.500 ;
    END
  END b10_not
  PIN a11_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 66.240 116.010 67.520 116.390 ;
        RECT 52.740 113.610 53.925 113.990 ;
        RECT 66.240 113.610 67.255 113.990 ;
        RECT 10.080 112.450 23.645 112.765 ;
        RECT 25.535 112.450 39.360 112.750 ;
        RECT 41.035 110.930 67.265 111.320 ;
        RECT 11.310 109.795 15.440 110.095 ;
        RECT 17.815 109.745 22.315 110.055 ;
        RECT 26.770 109.795 30.900 110.095 ;
        RECT 33.275 109.745 37.775 110.055 ;
        RECT 52.720 108.110 54.080 108.490 ;
        RECT 66.220 108.110 67.400 108.490 ;
        RECT 66.220 106.110 67.295 106.490 ;
      LAYER Metal2 ;
        RECT 10.085 112.405 10.465 112.785 ;
        RECT 23.250 112.405 23.630 112.785 ;
        RECT 25.520 112.405 25.900 112.810 ;
        RECT 38.985 112.405 39.345 114.235 ;
        RECT 41.165 110.885 41.580 114.235 ;
        RECT 53.360 113.975 53.670 114.005 ;
        RECT 53.360 107.875 53.675 113.975 ;
        RECT 66.860 105.880 67.190 116.575 ;
      LAYER Metal3 ;
        RECT 38.930 113.850 41.635 114.190 ;
        RECT 7.675 112.445 10.500 112.750 ;
        RECT 23.195 112.435 25.940 112.765 ;
    END
  END a11_f
  PIN a11_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 42.545 115.910 44.000 116.290 ;
        RECT 42.705 113.610 44.000 113.990 ;
        RECT 56.190 113.610 57.500 113.990 ;
        RECT 41.035 112.285 57.045 112.660 ;
        RECT 10.075 111.705 23.635 112.005 ;
        RECT 25.540 111.705 43.960 112.005 ;
        RECT 12.540 108.030 15.460 108.330 ;
        RECT 19.005 108.015 22.375 108.315 ;
        RECT 28.000 108.030 30.920 108.330 ;
        RECT 34.465 108.015 37.835 108.315 ;
        RECT 42.715 108.110 44.020 108.490 ;
        RECT 56.055 108.110 57.520 108.490 ;
        RECT 42.530 106.110 44.020 106.490 ;
      LAYER Metal2 ;
        RECT 10.075 111.655 10.455 112.035 ;
        RECT 12.575 107.980 12.875 112.040 ;
        RECT 19.065 107.965 19.345 112.055 ;
        RECT 23.255 111.655 23.635 112.035 ;
        RECT 25.525 111.655 25.905 112.060 ;
        RECT 28.035 107.980 28.335 112.040 ;
        RECT 34.525 107.965 34.805 112.055 ;
        RECT 42.835 106.055 43.190 116.360 ;
        RECT 43.500 111.660 43.845 112.715 ;
        RECT 56.345 107.830 56.675 114.025 ;
      LAYER Metal3 ;
        RECT 7.635 111.710 10.480 112.005 ;
        RECT 23.200 111.685 25.940 112.015 ;
    END
  END a11_not_f
  PIN b11
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 17.225 113.675 17.605 114.055 ;
        RECT 15.625 113.160 16.825 113.450 ;
        RECT 10.095 110.990 16.820 111.290 ;
        RECT 16.415 107.385 17.605 107.670 ;
        RECT 15.635 106.720 16.015 107.100 ;
      LAYER Metal2 ;
        RECT 10.120 110.970 10.500 111.350 ;
        RECT 15.675 106.710 15.975 113.520 ;
        RECT 16.465 107.305 16.775 113.495 ;
        RECT 17.260 107.235 17.560 114.065 ;
      LAYER Metal3 ;
        RECT 7.640 110.995 10.515 111.290 ;
    END
  END b11
  PIN b11_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT 10.765 113.875 14.140 114.275 ;
        RECT 22.545 113.225 22.925 113.605 ;
        RECT 10.075 110.370 14.200 110.640 ;
        RECT 13.775 109.195 20.165 109.485 ;
        RECT 10.755 107.280 11.135 107.660 ;
        RECT 19.755 106.555 22.935 106.875 ;
      LAYER Metal2 ;
        RECT 10.085 110.300 10.465 110.680 ;
        RECT 10.800 107.225 11.100 114.265 ;
        RECT 13.825 109.095 14.145 114.255 ;
        RECT 19.835 106.495 20.115 109.530 ;
        RECT 22.585 106.450 22.885 113.605 ;
      LAYER Metal3 ;
        RECT 7.675 110.365 10.470 110.660 ;
    END
  END b11_not
  PIN a12_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 66.110 96.300 67.390 96.680 ;
        RECT 52.610 93.900 53.795 94.280 ;
        RECT 66.110 93.900 67.125 94.280 ;
        RECT 9.950 92.740 23.515 93.055 ;
        RECT 25.405 92.740 39.230 93.040 ;
        RECT 40.905 91.220 67.135 91.610 ;
        RECT 11.180 90.085 15.310 90.385 ;
        RECT 17.685 90.035 22.185 90.345 ;
        RECT 26.640 90.085 30.770 90.385 ;
        RECT 33.145 90.035 37.645 90.345 ;
        RECT 52.590 88.400 53.950 88.780 ;
        RECT 66.090 88.400 67.270 88.780 ;
        RECT 66.090 86.400 67.165 86.780 ;
      LAYER Metal2 ;
        RECT 9.955 92.695 10.335 93.075 ;
        RECT 23.120 92.695 23.500 93.075 ;
        RECT 25.390 92.695 25.770 93.100 ;
        RECT 38.855 92.695 39.215 94.525 ;
        RECT 41.035 91.175 41.450 94.525 ;
        RECT 53.230 94.265 53.540 94.295 ;
        RECT 53.230 88.165 53.545 94.265 ;
        RECT 66.730 86.170 67.060 96.865 ;
      LAYER Metal3 ;
        RECT 38.800 94.140 41.505 94.480 ;
        RECT 7.545 92.735 10.370 93.040 ;
        RECT 23.065 92.725 25.810 93.055 ;
    END
  END a12_f
  PIN a12_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 42.415 96.200 43.870 96.580 ;
        RECT 42.575 93.900 43.870 94.280 ;
        RECT 56.060 93.900 57.370 94.280 ;
        RECT 40.905 92.575 56.915 92.950 ;
        RECT 9.945 91.995 23.505 92.295 ;
        RECT 25.410 91.995 43.830 92.295 ;
        RECT 12.410 88.320 15.330 88.620 ;
        RECT 18.875 88.305 22.245 88.605 ;
        RECT 27.870 88.320 30.790 88.620 ;
        RECT 34.335 88.305 37.705 88.605 ;
        RECT 42.585 88.400 43.890 88.780 ;
        RECT 55.925 88.400 57.390 88.780 ;
        RECT 42.400 86.400 43.890 86.780 ;
      LAYER Metal2 ;
        RECT 9.945 91.945 10.325 92.325 ;
        RECT 12.445 88.270 12.745 92.330 ;
        RECT 18.935 88.255 19.215 92.345 ;
        RECT 23.125 91.945 23.505 92.325 ;
        RECT 25.395 91.945 25.775 92.350 ;
        RECT 27.905 88.270 28.205 92.330 ;
        RECT 34.395 88.255 34.675 92.345 ;
        RECT 42.705 86.345 43.060 96.650 ;
        RECT 43.370 91.950 43.715 93.005 ;
        RECT 56.215 88.120 56.545 94.315 ;
      LAYER Metal3 ;
        RECT 7.505 92.000 10.350 92.295 ;
        RECT 23.070 91.975 25.810 92.305 ;
    END
  END a12_not_f
  PIN b12
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 17.095 93.965 17.475 94.345 ;
        RECT 15.495 93.450 16.695 93.740 ;
        RECT 9.965 91.280 16.690 91.580 ;
        RECT 16.285 87.675 17.475 87.960 ;
        RECT 15.505 87.010 15.885 87.390 ;
      LAYER Metal2 ;
        RECT 9.990 91.260 10.370 91.640 ;
        RECT 15.545 87.000 15.845 93.810 ;
        RECT 16.335 87.595 16.645 93.785 ;
        RECT 17.130 87.525 17.430 94.355 ;
      LAYER Metal3 ;
        RECT 7.510 91.285 10.385 91.580 ;
    END
  END b12
  PIN a8_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 102.905 175.195 104.140 175.575 ;
        RECT 100.880 172.795 104.140 173.175 ;
        RECT 108.310 171.635 121.925 171.935 ;
        RECT 109.505 168.980 113.635 169.280 ;
        RECT 116.010 168.930 120.510 169.240 ;
        RECT 102.765 167.935 106.710 168.270 ;
        RECT 100.860 167.295 104.160 167.675 ;
        RECT 102.675 165.295 104.160 165.675 ;
      LAYER Metal2 ;
        RECT 102.990 165.050 103.305 175.735 ;
        RECT 106.315 167.920 106.695 168.300 ;
        RECT 108.380 167.895 108.690 172.015 ;
        RECT 121.450 171.590 121.745 176.960 ;
      LAYER Metal3 ;
        RECT 121.450 176.505 137.470 176.915 ;
        RECT 106.315 167.910 108.795 168.310 ;
    END
  END a8_b
  PIN a10_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 83.335 135.725 84.535 136.105 ;
        RECT 83.335 133.425 86.595 133.805 ;
        RECT 84.000 131.510 106.555 131.850 ;
        RECT 107.665 131.520 122.310 131.820 ;
        RECT 83.315 127.925 86.615 128.305 ;
        RECT 110.690 127.845 113.610 128.145 ;
        RECT 117.155 127.830 120.525 128.130 ;
        RECT 83.315 125.925 84.600 126.305 ;
      LAYER Metal2 ;
        RECT 84.160 125.195 84.475 136.245 ;
        RECT 106.135 131.440 106.555 131.900 ;
        RECT 107.635 131.435 108.055 131.895 ;
        RECT 110.725 127.795 111.025 131.855 ;
        RECT 117.215 127.780 117.495 131.870 ;
        RECT 121.980 131.390 122.285 136.865 ;
      LAYER Metal3 ;
        RECT 121.935 136.355 137.415 136.810 ;
        RECT 106.105 131.490 108.130 131.875 ;
    END
  END a10_not_b
  PIN a11_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 102.860 116.030 104.095 116.410 ;
        RECT 100.835 113.630 104.095 114.010 ;
        RECT 108.265 112.470 121.880 112.770 ;
        RECT 109.460 109.815 113.590 110.115 ;
        RECT 115.965 109.765 120.465 110.075 ;
        RECT 102.720 108.770 106.665 109.105 ;
        RECT 100.815 108.130 104.115 108.510 ;
        RECT 102.630 106.130 104.115 106.510 ;
      LAYER Metal2 ;
        RECT 102.945 105.885 103.260 116.570 ;
        RECT 106.270 108.755 106.650 109.135 ;
        RECT 108.335 108.730 108.645 112.850 ;
        RECT 121.405 112.425 121.700 117.795 ;
      LAYER Metal3 ;
        RECT 121.405 117.340 137.425 117.750 ;
        RECT 106.270 108.745 108.750 109.145 ;
    END
  END a11_b
  PIN a11_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 83.335 115.930 84.535 116.310 ;
        RECT 83.335 113.630 86.595 114.010 ;
        RECT 84.000 111.715 106.555 112.055 ;
        RECT 107.665 111.725 122.310 112.025 ;
        RECT 83.315 108.130 86.615 108.510 ;
        RECT 110.690 108.050 113.610 108.350 ;
        RECT 117.155 108.035 120.525 108.335 ;
        RECT 83.315 106.130 84.600 106.510 ;
      LAYER Metal2 ;
        RECT 84.160 105.400 84.475 116.450 ;
        RECT 106.135 111.645 106.555 112.105 ;
        RECT 107.635 111.640 108.055 112.100 ;
        RECT 110.725 108.000 111.025 112.060 ;
        RECT 117.215 107.985 117.495 112.075 ;
        RECT 121.980 111.595 122.285 117.070 ;
      LAYER Metal3 ;
        RECT 121.935 116.560 137.415 117.015 ;
        RECT 106.105 111.695 108.130 112.080 ;
    END
  END a11_not_b
  PIN a12_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 102.780 96.275 104.015 96.655 ;
        RECT 100.755 93.875 104.015 94.255 ;
        RECT 108.185 92.715 121.800 93.015 ;
        RECT 109.380 90.060 113.510 90.360 ;
        RECT 115.885 90.010 120.385 90.320 ;
        RECT 102.640 89.015 106.585 89.350 ;
        RECT 100.735 88.375 104.035 88.755 ;
        RECT 102.550 86.375 104.035 86.755 ;
      LAYER Metal2 ;
        RECT 102.865 86.130 103.180 96.815 ;
        RECT 106.190 89.000 106.570 89.380 ;
        RECT 108.255 88.975 108.565 93.095 ;
        RECT 121.325 92.670 121.620 98.040 ;
      LAYER Metal3 ;
        RECT 121.325 97.585 137.345 97.995 ;
        RECT 106.190 88.990 108.670 89.390 ;
    END
  END a12_b
  PIN a12_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 83.255 96.175 84.455 96.555 ;
        RECT 83.255 93.875 86.515 94.255 ;
        RECT 83.920 91.960 106.475 92.300 ;
        RECT 107.585 91.970 122.230 92.270 ;
        RECT 83.235 88.375 86.535 88.755 ;
        RECT 110.610 88.295 113.530 88.595 ;
        RECT 117.075 88.280 120.445 88.580 ;
        RECT 83.235 86.375 84.520 86.755 ;
      LAYER Metal2 ;
        RECT 84.080 85.645 84.395 96.695 ;
        RECT 106.055 91.890 106.475 92.350 ;
        RECT 107.555 91.885 107.975 92.345 ;
        RECT 110.645 88.245 110.945 92.305 ;
        RECT 117.135 88.230 117.415 92.320 ;
        RECT 121.900 91.840 122.205 97.315 ;
      LAYER Metal3 ;
        RECT 121.855 96.805 137.335 97.260 ;
        RECT 106.025 91.940 108.050 92.325 ;
    END
  END a12_not_b
  PIN a13_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 102.885 76.560 104.120 76.940 ;
        RECT 100.860 74.160 104.120 74.540 ;
        RECT 108.290 73.000 121.905 73.300 ;
        RECT 109.485 70.345 113.615 70.645 ;
        RECT 115.990 70.295 120.490 70.605 ;
        RECT 102.745 69.300 106.690 69.635 ;
        RECT 100.840 68.660 104.140 69.040 ;
        RECT 102.655 66.660 104.140 67.040 ;
      LAYER Metal2 ;
        RECT 102.970 66.415 103.285 77.100 ;
        RECT 106.295 69.285 106.675 69.665 ;
        RECT 108.360 69.260 108.670 73.380 ;
        RECT 121.430 72.955 121.725 78.325 ;
      LAYER Metal3 ;
        RECT 121.430 77.870 137.450 78.280 ;
        RECT 106.295 69.275 108.775 69.675 ;
    END
  END a13_b
  PIN a13_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 83.360 76.460 84.560 76.840 ;
        RECT 83.360 74.160 86.620 74.540 ;
        RECT 84.025 72.245 106.580 72.585 ;
        RECT 107.690 72.255 122.335 72.555 ;
        RECT 83.340 68.660 86.640 69.040 ;
        RECT 110.715 68.580 113.635 68.880 ;
        RECT 117.180 68.565 120.550 68.865 ;
        RECT 83.340 66.660 84.625 67.040 ;
      LAYER Metal2 ;
        RECT 84.185 65.930 84.500 76.980 ;
        RECT 106.160 72.175 106.580 72.635 ;
        RECT 107.660 72.170 108.080 72.630 ;
        RECT 110.750 68.530 111.050 72.590 ;
        RECT 117.240 68.515 117.520 72.605 ;
        RECT 122.005 72.125 122.310 77.600 ;
      LAYER Metal3 ;
        RECT 121.960 77.090 137.440 77.545 ;
        RECT 106.130 72.225 108.155 72.610 ;
    END
  END a13_not_b
  PIN a14_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 102.885 56.590 104.120 56.970 ;
        RECT 100.860 54.190 104.120 54.570 ;
        RECT 108.290 53.030 121.905 53.330 ;
        RECT 109.485 50.375 113.615 50.675 ;
        RECT 115.990 50.325 120.490 50.635 ;
        RECT 102.745 49.330 106.690 49.665 ;
        RECT 100.840 48.690 104.140 49.070 ;
        RECT 102.655 46.690 104.140 47.070 ;
      LAYER Metal2 ;
        RECT 102.970 46.445 103.285 57.130 ;
        RECT 106.295 49.315 106.675 49.695 ;
        RECT 108.360 49.290 108.670 53.410 ;
        RECT 121.430 52.985 121.725 58.355 ;
      LAYER Metal3 ;
        RECT 121.430 57.900 137.450 58.310 ;
        RECT 106.295 49.305 108.775 49.705 ;
    END
  END a14_b
  PIN a14_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 83.360 56.490 84.560 56.870 ;
        RECT 83.360 54.190 86.620 54.570 ;
        RECT 84.025 52.275 106.580 52.615 ;
        RECT 107.690 52.285 122.335 52.585 ;
        RECT 83.340 48.690 86.640 49.070 ;
        RECT 110.715 48.610 113.635 48.910 ;
        RECT 117.180 48.595 120.550 48.895 ;
        RECT 83.340 46.690 84.625 47.070 ;
      LAYER Metal2 ;
        RECT 84.185 45.960 84.500 57.010 ;
        RECT 106.160 52.205 106.580 52.665 ;
        RECT 107.660 52.200 108.080 52.660 ;
        RECT 110.750 48.560 111.050 52.620 ;
        RECT 117.240 48.545 117.520 52.635 ;
        RECT 122.005 52.155 122.310 57.630 ;
      LAYER Metal3 ;
        RECT 121.960 57.120 137.440 57.575 ;
        RECT 106.130 52.255 108.155 52.640 ;
    END
  END a14_not_b
  PIN a15_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 102.885 36.925 104.120 37.305 ;
        RECT 100.860 34.525 104.120 34.905 ;
        RECT 108.290 33.365 121.905 33.665 ;
        RECT 109.485 30.710 113.615 31.010 ;
        RECT 115.990 30.660 120.490 30.970 ;
        RECT 102.745 29.665 106.690 30.000 ;
        RECT 100.840 29.025 104.140 29.405 ;
        RECT 102.655 27.025 104.140 27.405 ;
      LAYER Metal2 ;
        RECT 102.970 26.780 103.285 37.465 ;
        RECT 106.295 29.650 106.675 30.030 ;
        RECT 108.360 29.625 108.670 33.745 ;
        RECT 121.430 33.320 121.725 38.690 ;
      LAYER Metal3 ;
        RECT 121.430 38.235 137.450 38.645 ;
        RECT 106.295 29.640 108.775 30.040 ;
    END
  END a15_b
  PIN a15_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 83.360 36.825 84.560 37.205 ;
        RECT 83.360 34.525 86.620 34.905 ;
        RECT 84.025 32.610 106.580 32.950 ;
        RECT 107.690 32.620 122.335 32.920 ;
        RECT 83.340 29.025 86.640 29.405 ;
        RECT 110.715 28.945 113.635 29.245 ;
        RECT 117.180 28.930 120.550 29.230 ;
        RECT 83.340 27.025 84.625 27.405 ;
      LAYER Metal2 ;
        RECT 84.185 26.295 84.500 37.345 ;
        RECT 106.160 32.540 106.580 33.000 ;
        RECT 107.660 32.535 108.080 32.995 ;
        RECT 110.750 28.895 111.050 32.955 ;
        RECT 117.240 28.880 117.520 32.970 ;
        RECT 122.005 32.490 122.310 37.965 ;
      LAYER Metal3 ;
        RECT 121.960 37.455 137.440 37.910 ;
        RECT 106.130 32.590 108.155 32.975 ;
    END
  END a15_not_b
  PIN a8_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 83.380 175.095 84.580 175.475 ;
        RECT 83.380 172.795 86.640 173.175 ;
        RECT 84.045 170.880 106.600 171.220 ;
        RECT 107.710 170.890 122.355 171.190 ;
        RECT 83.360 167.295 86.660 167.675 ;
        RECT 110.735 167.215 113.655 167.515 ;
        RECT 117.200 167.200 120.570 167.500 ;
        RECT 83.360 165.295 84.645 165.675 ;
      LAYER Metal2 ;
        RECT 84.205 164.565 84.520 175.615 ;
        RECT 106.180 170.810 106.600 171.270 ;
        RECT 107.680 170.805 108.100 171.265 ;
        RECT 110.770 167.165 111.070 171.225 ;
        RECT 117.260 167.150 117.540 171.240 ;
        RECT 122.025 170.760 122.330 176.235 ;
      LAYER Metal3 ;
        RECT 121.980 175.725 137.460 176.180 ;
        RECT 106.150 170.860 108.175 171.245 ;
    END
  END a8_not_b
  PIN a9_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 102.705 155.470 103.940 155.850 ;
        RECT 100.680 153.070 103.940 153.450 ;
        RECT 108.110 151.910 121.725 152.210 ;
        RECT 109.305 149.255 113.435 149.555 ;
        RECT 115.810 149.205 120.310 149.515 ;
        RECT 102.565 148.210 106.510 148.545 ;
        RECT 100.660 147.570 103.960 147.950 ;
        RECT 102.475 145.570 103.960 145.950 ;
      LAYER Metal2 ;
        RECT 102.790 145.325 103.105 156.010 ;
        RECT 106.115 148.195 106.495 148.575 ;
        RECT 108.180 148.170 108.490 152.290 ;
        RECT 121.250 151.865 121.545 157.235 ;
      LAYER Metal3 ;
        RECT 121.250 156.780 137.270 157.190 ;
        RECT 106.115 148.185 108.595 148.585 ;
    END
  END a9_b
  PIN a9_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 83.180 155.370 84.380 155.750 ;
        RECT 83.180 153.070 86.440 153.450 ;
        RECT 83.845 151.155 106.400 151.495 ;
        RECT 107.510 151.165 122.155 151.465 ;
        RECT 83.160 147.570 86.460 147.950 ;
        RECT 110.535 147.490 113.455 147.790 ;
        RECT 117.000 147.475 120.370 147.775 ;
        RECT 83.160 145.570 84.445 145.950 ;
      LAYER Metal2 ;
        RECT 84.005 144.840 84.320 155.890 ;
        RECT 105.980 151.085 106.400 151.545 ;
        RECT 107.480 151.080 107.900 151.540 ;
        RECT 110.570 147.440 110.870 151.500 ;
        RECT 117.060 147.425 117.340 151.515 ;
        RECT 121.825 151.035 122.130 156.510 ;
      LAYER Metal3 ;
        RECT 121.780 156.000 137.260 156.455 ;
        RECT 105.950 151.135 107.975 151.520 ;
    END
  END a9_not_b
  PIN a10_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 102.860 135.825 104.095 136.205 ;
        RECT 100.835 133.425 104.095 133.805 ;
        RECT 108.265 132.265 121.880 132.565 ;
        RECT 109.460 129.610 113.590 129.910 ;
        RECT 115.965 129.560 120.465 129.870 ;
        RECT 102.720 128.565 106.665 128.900 ;
        RECT 100.815 127.925 104.115 128.305 ;
        RECT 102.630 125.925 104.115 126.305 ;
      LAYER Metal2 ;
        RECT 102.945 125.680 103.260 136.365 ;
        RECT 106.270 128.550 106.650 128.930 ;
        RECT 108.335 128.525 108.645 132.645 ;
        RECT 121.405 132.220 121.700 137.590 ;
      LAYER Metal3 ;
        RECT 121.405 137.135 137.425 137.545 ;
        RECT 106.270 128.540 108.750 128.940 ;
    END
  END a10_b
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 8.165 320.415 39.085 328.115 ;
        RECT 41.065 320.415 67.720 328.115 ;
        RECT 79.655 320.360 137.230 328.060 ;
        RECT 8.120 300.725 39.040 308.425 ;
        RECT 41.020 300.725 67.675 308.425 ;
        RECT 79.455 300.635 137.030 308.335 ;
        RECT 8.310 281.015 39.230 288.715 ;
        RECT 41.210 281.015 67.865 288.715 ;
        RECT 79.610 280.990 137.185 288.690 ;
        RECT 8.115 261.175 39.035 268.875 ;
        RECT 41.015 261.175 67.670 268.875 ;
        RECT 79.610 261.195 137.185 268.895 ;
        RECT 7.985 241.465 38.905 249.165 ;
        RECT 40.885 241.465 67.540 249.165 ;
        RECT 79.530 241.440 137.105 249.140 ;
        RECT 8.115 221.705 39.035 229.405 ;
        RECT 41.015 221.705 67.670 229.405 ;
        RECT 79.635 221.725 137.210 229.425 ;
        RECT 8.065 201.895 38.985 209.595 ;
        RECT 40.965 201.895 67.620 209.595 ;
        RECT 79.635 201.755 137.210 209.455 ;
        RECT 8.035 182.100 38.955 189.800 ;
        RECT 40.935 182.100 67.590 189.800 ;
        RECT 79.635 182.090 137.210 189.790 ;
        RECT 8.185 162.305 39.105 170.005 ;
        RECT 41.085 162.305 67.740 170.005 ;
        RECT 79.675 162.250 137.250 169.950 ;
        RECT 8.140 142.615 39.060 150.315 ;
        RECT 41.040 142.615 67.695 150.315 ;
        RECT 79.475 142.525 137.050 150.225 ;
        RECT 8.330 122.905 39.250 130.605 ;
        RECT 41.230 122.905 67.885 130.605 ;
        RECT 79.630 122.880 137.205 130.580 ;
        RECT 8.135 103.065 39.055 110.765 ;
        RECT 41.035 103.065 67.690 110.765 ;
        RECT 79.630 103.085 137.205 110.785 ;
        RECT 8.005 83.355 38.925 91.055 ;
        RECT 40.905 83.355 67.560 91.055 ;
        RECT 79.550 83.330 137.125 91.030 ;
        RECT 8.135 63.595 39.055 71.295 ;
        RECT 41.035 63.595 67.690 71.295 ;
        RECT 79.655 63.615 137.230 71.315 ;
        RECT 8.085 43.785 39.005 51.485 ;
        RECT 40.985 43.785 67.640 51.485 ;
        RECT 79.655 43.645 137.230 51.345 ;
        RECT 8.055 23.990 38.975 31.690 ;
        RECT 40.955 23.990 67.610 31.690 ;
        RECT 79.655 23.980 137.230 31.680 ;
        RECT 79.670 4.245 95.130 11.945 ;
      LAYER Metal1 ;
        RECT 8.965 321.315 9.345 327.145 ;
        RECT 9.715 321.315 13.810 321.320 ;
        RECT 24.425 321.315 24.805 327.145 ;
        RECT 46.255 322.780 47.775 323.140 ;
        RECT 84.845 322.725 86.365 323.085 ;
        RECT 25.175 321.315 29.270 321.320 ;
        RECT 8.595 321.310 13.810 321.315 ;
        RECT 24.055 321.310 29.270 321.315 ;
        RECT 39.515 321.310 79.765 321.315 ;
        RECT 8.595 321.260 79.765 321.310 ;
        RECT 106.310 321.260 111.955 321.265 ;
        RECT 122.570 321.260 122.950 327.090 ;
        RECT 123.320 321.260 127.415 321.265 ;
        RECT 8.595 321.255 111.955 321.260 ;
        RECT 122.200 321.255 127.415 321.260 ;
        RECT 8.595 320.415 137.230 321.255 ;
        RECT 79.655 320.360 137.230 320.415 ;
        RECT 8.920 301.625 9.300 307.455 ;
        RECT 9.670 301.625 13.765 301.630 ;
        RECT 24.380 301.625 24.760 307.455 ;
        RECT 46.210 303.090 47.730 303.450 ;
        RECT 84.645 303.000 86.165 303.360 ;
        RECT 25.130 301.625 29.225 301.630 ;
        RECT 8.550 301.620 13.765 301.625 ;
        RECT 24.010 301.620 29.225 301.625 ;
        RECT 39.470 301.620 79.720 301.625 ;
        RECT 8.550 301.535 79.720 301.620 ;
        RECT 106.110 301.535 111.755 301.540 ;
        RECT 122.370 301.535 122.750 307.365 ;
        RECT 123.120 301.535 127.215 301.540 ;
        RECT 8.550 301.530 111.755 301.535 ;
        RECT 122.000 301.530 127.215 301.535 ;
        RECT 8.550 300.725 137.030 301.530 ;
        RECT 79.455 300.635 137.030 300.725 ;
        RECT 9.110 281.915 9.490 287.745 ;
        RECT 9.860 281.915 13.955 281.920 ;
        RECT 24.570 281.915 24.950 287.745 ;
        RECT 46.400 283.380 47.920 283.740 ;
        RECT 84.800 283.355 86.320 283.715 ;
        RECT 25.320 281.915 29.415 281.920 ;
        RECT 8.740 281.910 13.955 281.915 ;
        RECT 24.200 281.910 29.415 281.915 ;
        RECT 39.660 281.910 79.910 281.915 ;
        RECT 8.740 281.890 79.910 281.910 ;
        RECT 106.265 281.890 111.910 281.895 ;
        RECT 122.525 281.890 122.905 287.720 ;
        RECT 123.275 281.890 127.370 281.895 ;
        RECT 8.740 281.885 111.910 281.890 ;
        RECT 122.155 281.885 127.370 281.890 ;
        RECT 8.740 281.015 137.185 281.885 ;
        RECT 79.610 280.990 137.185 281.015 ;
        RECT 8.915 262.075 9.295 267.905 ;
        RECT 9.665 262.075 13.760 262.080 ;
        RECT 24.375 262.075 24.755 267.905 ;
        RECT 46.205 263.540 47.725 263.900 ;
        RECT 84.800 263.560 86.320 263.920 ;
        RECT 106.265 262.095 111.910 262.100 ;
        RECT 122.525 262.095 122.905 267.925 ;
        RECT 123.275 262.095 127.370 262.100 ;
        RECT 79.610 262.090 111.910 262.095 ;
        RECT 122.155 262.090 127.370 262.095 ;
        RECT 25.125 262.075 29.220 262.080 ;
        RECT 79.610 262.075 137.185 262.090 ;
        RECT 8.545 262.070 13.760 262.075 ;
        RECT 24.005 262.070 29.220 262.075 ;
        RECT 39.465 262.070 137.185 262.075 ;
        RECT 8.545 261.195 137.185 262.070 ;
        RECT 8.545 261.175 79.715 261.195 ;
        RECT 8.785 242.365 9.165 248.195 ;
        RECT 9.535 242.365 13.630 242.370 ;
        RECT 24.245 242.365 24.625 248.195 ;
        RECT 46.075 243.830 47.595 244.190 ;
        RECT 84.720 243.805 86.240 244.165 ;
        RECT 24.995 242.365 29.090 242.370 ;
        RECT 8.415 242.360 13.630 242.365 ;
        RECT 23.875 242.360 29.090 242.365 ;
        RECT 39.335 242.360 79.585 242.365 ;
        RECT 8.415 242.340 79.585 242.360 ;
        RECT 106.185 242.340 111.830 242.345 ;
        RECT 122.445 242.340 122.825 248.170 ;
        RECT 123.195 242.340 127.290 242.345 ;
        RECT 8.415 242.335 111.830 242.340 ;
        RECT 122.075 242.335 127.290 242.340 ;
        RECT 8.415 241.465 137.105 242.335 ;
        RECT 79.530 241.440 137.105 241.465 ;
        RECT 8.915 222.605 9.295 228.435 ;
        RECT 9.665 222.605 13.760 222.610 ;
        RECT 24.375 222.605 24.755 228.435 ;
        RECT 46.205 224.070 47.725 224.430 ;
        RECT 84.825 224.090 86.345 224.450 ;
        RECT 106.290 222.625 111.935 222.630 ;
        RECT 122.550 222.625 122.930 228.455 ;
        RECT 123.300 222.625 127.395 222.630 ;
        RECT 79.635 222.620 111.935 222.625 ;
        RECT 122.180 222.620 127.395 222.625 ;
        RECT 25.125 222.605 29.220 222.610 ;
        RECT 79.635 222.605 137.210 222.620 ;
        RECT 8.545 222.600 13.760 222.605 ;
        RECT 24.005 222.600 29.220 222.605 ;
        RECT 39.465 222.600 137.210 222.605 ;
        RECT 8.545 221.725 137.210 222.600 ;
        RECT 8.545 221.705 79.715 221.725 ;
        RECT 8.865 202.795 9.245 208.625 ;
        RECT 9.615 202.795 13.710 202.800 ;
        RECT 24.325 202.795 24.705 208.625 ;
        RECT 46.155 204.260 47.675 204.620 ;
        RECT 84.825 204.120 86.345 204.480 ;
        RECT 25.075 202.795 29.170 202.800 ;
        RECT 8.495 202.790 13.710 202.795 ;
        RECT 23.955 202.790 29.170 202.795 ;
        RECT 39.415 202.790 79.665 202.795 ;
        RECT 8.495 202.655 79.665 202.790 ;
        RECT 106.290 202.655 111.935 202.660 ;
        RECT 122.550 202.655 122.930 208.485 ;
        RECT 123.300 202.655 127.395 202.660 ;
        RECT 8.495 202.650 111.935 202.655 ;
        RECT 122.180 202.650 127.395 202.655 ;
        RECT 8.495 201.895 137.210 202.650 ;
        RECT 79.635 201.755 137.210 201.895 ;
        RECT 8.835 183.000 9.215 188.830 ;
        RECT 9.585 183.000 13.680 183.005 ;
        RECT 24.295 183.000 24.675 188.830 ;
        RECT 46.125 184.465 47.645 184.825 ;
        RECT 84.825 184.455 86.345 184.815 ;
        RECT 25.045 183.000 29.140 183.005 ;
        RECT 8.465 182.995 13.680 183.000 ;
        RECT 23.925 182.995 29.140 183.000 ;
        RECT 39.385 182.995 79.635 183.000 ;
        RECT 8.465 182.990 79.635 182.995 ;
        RECT 106.290 182.990 111.935 182.995 ;
        RECT 122.550 182.990 122.930 188.820 ;
        RECT 123.300 182.990 127.395 182.995 ;
        RECT 8.465 182.985 111.935 182.990 ;
        RECT 122.180 182.985 127.395 182.990 ;
        RECT 8.465 182.100 137.210 182.985 ;
        RECT 79.635 182.090 137.210 182.100 ;
        RECT 8.985 163.205 9.365 169.035 ;
        RECT 9.735 163.205 13.830 163.210 ;
        RECT 24.445 163.205 24.825 169.035 ;
        RECT 46.275 164.670 47.795 165.030 ;
        RECT 84.865 164.615 86.385 164.975 ;
        RECT 25.195 163.205 29.290 163.210 ;
        RECT 8.615 163.200 13.830 163.205 ;
        RECT 24.075 163.200 29.290 163.205 ;
        RECT 39.535 163.200 79.785 163.205 ;
        RECT 8.615 163.150 79.785 163.200 ;
        RECT 106.330 163.150 111.975 163.155 ;
        RECT 122.590 163.150 122.970 168.980 ;
        RECT 123.340 163.150 127.435 163.155 ;
        RECT 8.615 163.145 111.975 163.150 ;
        RECT 122.220 163.145 127.435 163.150 ;
        RECT 8.615 162.305 137.250 163.145 ;
        RECT 79.675 162.250 137.250 162.305 ;
        RECT 8.940 143.515 9.320 149.345 ;
        RECT 9.690 143.515 13.785 143.520 ;
        RECT 24.400 143.515 24.780 149.345 ;
        RECT 46.230 144.980 47.750 145.340 ;
        RECT 84.665 144.890 86.185 145.250 ;
        RECT 25.150 143.515 29.245 143.520 ;
        RECT 8.570 143.510 13.785 143.515 ;
        RECT 24.030 143.510 29.245 143.515 ;
        RECT 39.490 143.510 79.740 143.515 ;
        RECT 8.570 143.425 79.740 143.510 ;
        RECT 106.130 143.425 111.775 143.430 ;
        RECT 122.390 143.425 122.770 149.255 ;
        RECT 123.140 143.425 127.235 143.430 ;
        RECT 8.570 143.420 111.775 143.425 ;
        RECT 122.020 143.420 127.235 143.425 ;
        RECT 8.570 142.615 137.050 143.420 ;
        RECT 79.475 142.525 137.050 142.615 ;
        RECT 9.130 123.805 9.510 129.635 ;
        RECT 9.880 123.805 13.975 123.810 ;
        RECT 24.590 123.805 24.970 129.635 ;
        RECT 46.420 125.270 47.940 125.630 ;
        RECT 84.820 125.245 86.340 125.605 ;
        RECT 25.340 123.805 29.435 123.810 ;
        RECT 8.760 123.800 13.975 123.805 ;
        RECT 24.220 123.800 29.435 123.805 ;
        RECT 39.680 123.800 79.930 123.805 ;
        RECT 8.760 123.780 79.930 123.800 ;
        RECT 106.285 123.780 111.930 123.785 ;
        RECT 122.545 123.780 122.925 129.610 ;
        RECT 123.295 123.780 127.390 123.785 ;
        RECT 8.760 123.775 111.930 123.780 ;
        RECT 122.175 123.775 127.390 123.780 ;
        RECT 8.760 122.905 137.205 123.775 ;
        RECT 79.630 122.880 137.205 122.905 ;
        RECT 8.935 103.965 9.315 109.795 ;
        RECT 9.685 103.965 13.780 103.970 ;
        RECT 24.395 103.965 24.775 109.795 ;
        RECT 46.225 105.430 47.745 105.790 ;
        RECT 84.820 105.450 86.340 105.810 ;
        RECT 106.285 103.985 111.930 103.990 ;
        RECT 122.545 103.985 122.925 109.815 ;
        RECT 123.295 103.985 127.390 103.990 ;
        RECT 79.630 103.980 111.930 103.985 ;
        RECT 122.175 103.980 127.390 103.985 ;
        RECT 25.145 103.965 29.240 103.970 ;
        RECT 79.630 103.965 137.205 103.980 ;
        RECT 8.565 103.960 13.780 103.965 ;
        RECT 24.025 103.960 29.240 103.965 ;
        RECT 39.485 103.960 137.205 103.965 ;
        RECT 8.565 103.085 137.205 103.960 ;
        RECT 8.565 103.065 79.735 103.085 ;
        RECT 8.805 84.255 9.185 90.085 ;
        RECT 9.555 84.255 13.650 84.260 ;
        RECT 24.265 84.255 24.645 90.085 ;
        RECT 46.095 85.720 47.615 86.080 ;
        RECT 84.740 85.695 86.260 86.055 ;
        RECT 25.015 84.255 29.110 84.260 ;
        RECT 8.435 84.250 13.650 84.255 ;
        RECT 23.895 84.250 29.110 84.255 ;
        RECT 39.355 84.250 79.605 84.255 ;
        RECT 8.435 84.230 79.605 84.250 ;
        RECT 106.205 84.230 111.850 84.235 ;
        RECT 122.465 84.230 122.845 90.060 ;
        RECT 123.215 84.230 127.310 84.235 ;
        RECT 8.435 84.225 111.850 84.230 ;
        RECT 122.095 84.225 127.310 84.230 ;
        RECT 8.435 83.355 137.125 84.225 ;
        RECT 79.550 83.330 137.125 83.355 ;
        RECT 8.935 64.495 9.315 70.325 ;
        RECT 9.685 64.495 13.780 64.500 ;
        RECT 24.395 64.495 24.775 70.325 ;
        RECT 46.225 65.960 47.745 66.320 ;
        RECT 84.845 65.980 86.365 66.340 ;
        RECT 106.310 64.515 111.955 64.520 ;
        RECT 122.570 64.515 122.950 70.345 ;
        RECT 123.320 64.515 127.415 64.520 ;
        RECT 79.655 64.510 111.955 64.515 ;
        RECT 122.200 64.510 127.415 64.515 ;
        RECT 25.145 64.495 29.240 64.500 ;
        RECT 79.655 64.495 137.230 64.510 ;
        RECT 8.565 64.490 13.780 64.495 ;
        RECT 24.025 64.490 29.240 64.495 ;
        RECT 39.485 64.490 137.230 64.495 ;
        RECT 8.565 63.615 137.230 64.490 ;
        RECT 8.565 63.595 79.735 63.615 ;
        RECT 8.885 44.685 9.265 50.515 ;
        RECT 9.635 44.685 13.730 44.690 ;
        RECT 24.345 44.685 24.725 50.515 ;
        RECT 46.175 46.150 47.695 46.510 ;
        RECT 84.845 46.010 86.365 46.370 ;
        RECT 25.095 44.685 29.190 44.690 ;
        RECT 8.515 44.680 13.730 44.685 ;
        RECT 23.975 44.680 29.190 44.685 ;
        RECT 39.435 44.680 79.685 44.685 ;
        RECT 8.515 44.545 79.685 44.680 ;
        RECT 106.310 44.545 111.955 44.550 ;
        RECT 122.570 44.545 122.950 50.375 ;
        RECT 123.320 44.545 127.415 44.550 ;
        RECT 8.515 44.540 111.955 44.545 ;
        RECT 122.200 44.540 127.415 44.545 ;
        RECT 8.515 43.785 137.230 44.540 ;
        RECT 79.655 43.645 137.230 43.785 ;
        RECT 8.855 24.890 9.235 30.720 ;
        RECT 9.605 24.890 13.700 24.895 ;
        RECT 24.315 24.890 24.695 30.720 ;
        RECT 46.145 26.355 47.665 26.715 ;
        RECT 84.845 26.345 86.365 26.705 ;
        RECT 25.065 24.890 29.160 24.895 ;
        RECT 8.485 24.885 13.700 24.890 ;
        RECT 23.945 24.885 29.160 24.890 ;
        RECT 39.405 24.885 79.655 24.890 ;
        RECT 8.485 24.880 79.655 24.885 ;
        RECT 106.310 24.880 111.955 24.885 ;
        RECT 122.570 24.880 122.950 30.710 ;
        RECT 123.320 24.880 127.415 24.885 ;
        RECT 8.485 24.875 111.955 24.880 ;
        RECT 122.200 24.875 127.415 24.880 ;
        RECT 8.485 23.990 137.230 24.875 ;
        RECT 79.655 23.980 137.230 23.990 ;
        RECT 70.800 5.140 83.335 5.150 ;
        RECT 93.950 5.145 94.330 10.975 ;
        RECT 93.580 5.140 94.700 5.145 ;
        RECT 70.800 4.245 94.700 5.140 ;
      LAYER Metal2 ;
        RECT 47.265 320.880 47.610 323.340 ;
        RECT 47.220 301.190 47.565 303.650 ;
        RECT 47.410 281.480 47.755 283.940 ;
        RECT 47.215 261.640 47.560 264.100 ;
        RECT 47.085 241.930 47.430 244.390 ;
        RECT 47.215 222.170 47.560 224.630 ;
        RECT 47.165 202.360 47.510 204.820 ;
        RECT 47.135 182.565 47.480 185.025 ;
        RECT 47.285 162.770 47.630 165.230 ;
        RECT 47.240 143.080 47.585 145.540 ;
        RECT 47.430 123.370 47.775 125.830 ;
        RECT 47.235 103.530 47.580 105.990 ;
        RECT 47.105 83.820 47.450 86.280 ;
        RECT 47.235 64.060 47.580 66.520 ;
        RECT 47.185 44.250 47.530 46.710 ;
        RECT 47.155 24.455 47.500 26.915 ;
        RECT 70.800 4.195 71.215 336.340 ;
        RECT 85.855 320.825 86.200 323.285 ;
        RECT 85.655 301.100 86.000 303.560 ;
        RECT 85.810 281.455 86.155 283.915 ;
        RECT 85.810 261.660 86.155 264.120 ;
        RECT 85.730 241.905 86.075 244.365 ;
        RECT 85.835 222.190 86.180 224.650 ;
        RECT 85.835 202.220 86.180 204.680 ;
        RECT 85.835 182.555 86.180 185.015 ;
        RECT 85.875 162.715 86.220 165.175 ;
        RECT 85.675 142.990 86.020 145.450 ;
        RECT 85.830 123.345 86.175 125.805 ;
        RECT 85.830 103.550 86.175 106.010 ;
        RECT 85.750 83.795 86.095 86.255 ;
        RECT 85.855 64.080 86.200 66.540 ;
        RECT 85.855 44.110 86.200 46.570 ;
        RECT 85.855 24.445 86.200 26.905 ;
      LAYER Metal3 ;
        RECT 54.420 17.980 71.210 18.470 ;
      LAYER Metal4 ;
        RECT 59.520 13.840 60.765 18.470 ;
        RECT 54.565 2.790 65.770 13.840 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT 8.165 328.115 67.720 336.340 ;
        RECT 79.655 328.060 137.230 336.285 ;
        RECT 8.120 308.425 67.675 316.650 ;
        RECT 79.455 308.335 137.030 316.560 ;
        RECT 8.310 288.715 67.865 296.940 ;
        RECT 79.610 288.690 137.185 296.915 ;
        RECT 8.115 268.875 67.670 277.100 ;
        RECT 79.610 268.895 137.185 277.120 ;
        RECT 7.985 249.165 67.540 257.390 ;
        RECT 79.530 249.140 137.105 257.365 ;
        RECT 8.115 229.405 67.670 237.630 ;
        RECT 79.635 229.425 137.210 237.650 ;
        RECT 8.065 209.595 67.620 217.820 ;
        RECT 79.635 209.455 137.210 217.680 ;
        RECT 8.035 189.800 67.590 198.025 ;
        RECT 79.635 189.790 137.210 198.015 ;
        RECT 8.185 170.005 67.740 178.230 ;
        RECT 79.675 169.950 137.250 178.175 ;
        RECT 8.140 150.315 67.695 158.540 ;
        RECT 79.475 150.225 137.050 158.450 ;
        RECT 8.330 130.605 67.885 138.830 ;
        RECT 79.630 130.580 137.205 138.805 ;
        RECT 8.135 110.765 67.690 118.990 ;
        RECT 79.630 110.785 137.205 119.010 ;
        RECT 8.005 91.055 67.560 99.280 ;
        RECT 79.550 91.030 137.125 99.255 ;
        RECT 8.135 71.295 67.690 79.520 ;
        RECT 79.655 71.315 137.230 79.540 ;
        RECT 8.085 51.485 67.640 59.710 ;
        RECT 79.655 51.345 137.230 59.570 ;
        RECT 8.055 31.690 67.610 39.915 ;
        RECT 79.655 31.680 137.230 39.905 ;
        RECT 79.670 11.945 95.130 20.170 ;
      LAYER Metal1 ;
        RECT 8.595 336.285 80.985 336.340 ;
        RECT 8.595 335.440 137.230 336.285 ;
        RECT 8.965 328.280 9.345 335.440 ;
        RECT 24.425 328.280 24.805 335.440 ;
        RECT 80.875 335.385 137.230 335.440 ;
        RECT 47.725 333.045 50.000 333.555 ;
        RECT 52.625 333.045 54.925 333.555 ;
        RECT 57.220 333.045 59.500 333.555 ;
        RECT 86.315 332.990 88.590 333.500 ;
        RECT 91.215 332.990 93.515 333.500 ;
        RECT 95.810 332.990 98.090 333.500 ;
        RECT 122.570 328.225 122.950 335.385 ;
        RECT 8.550 316.560 80.940 316.650 ;
        RECT 8.550 315.750 137.030 316.560 ;
        RECT 8.920 308.590 9.300 315.750 ;
        RECT 24.380 308.590 24.760 315.750 ;
        RECT 80.675 315.660 137.030 315.750 ;
        RECT 47.680 313.355 49.955 313.865 ;
        RECT 52.580 313.355 54.880 313.865 ;
        RECT 57.175 313.355 59.455 313.865 ;
        RECT 86.115 313.265 88.390 313.775 ;
        RECT 91.015 313.265 93.315 313.775 ;
        RECT 95.610 313.265 97.890 313.775 ;
        RECT 122.370 308.500 122.750 315.660 ;
        RECT 8.740 296.915 81.130 296.940 ;
        RECT 8.740 296.040 137.185 296.915 ;
        RECT 9.110 288.880 9.490 296.040 ;
        RECT 24.570 288.880 24.950 296.040 ;
        RECT 80.830 296.015 137.185 296.040 ;
        RECT 47.870 293.645 50.145 294.155 ;
        RECT 52.770 293.645 55.070 294.155 ;
        RECT 57.365 293.645 59.645 294.155 ;
        RECT 86.270 293.620 88.545 294.130 ;
        RECT 91.170 293.620 93.470 294.130 ;
        RECT 95.765 293.620 98.045 294.130 ;
        RECT 122.525 288.855 122.905 296.015 ;
        RECT 80.830 277.100 137.185 277.120 ;
        RECT 8.545 276.220 137.185 277.100 ;
        RECT 8.545 276.200 80.935 276.220 ;
        RECT 8.915 269.040 9.295 276.200 ;
        RECT 24.375 269.040 24.755 276.200 ;
        RECT 47.675 273.805 49.950 274.315 ;
        RECT 52.575 273.805 54.875 274.315 ;
        RECT 57.170 273.805 59.450 274.315 ;
        RECT 86.270 273.825 88.545 274.335 ;
        RECT 91.170 273.825 93.470 274.335 ;
        RECT 95.765 273.825 98.045 274.335 ;
        RECT 122.525 269.060 122.905 276.220 ;
        RECT 8.415 257.365 80.805 257.390 ;
        RECT 8.415 256.490 137.105 257.365 ;
        RECT 8.785 249.330 9.165 256.490 ;
        RECT 24.245 249.330 24.625 256.490 ;
        RECT 80.750 256.465 137.105 256.490 ;
        RECT 47.545 254.095 49.820 254.605 ;
        RECT 52.445 254.095 54.745 254.605 ;
        RECT 57.040 254.095 59.320 254.605 ;
        RECT 86.190 254.070 88.465 254.580 ;
        RECT 91.090 254.070 93.390 254.580 ;
        RECT 95.685 254.070 97.965 254.580 ;
        RECT 122.445 249.305 122.825 256.465 ;
        RECT 80.855 237.630 137.210 237.650 ;
        RECT 8.545 236.750 137.210 237.630 ;
        RECT 8.545 236.730 80.935 236.750 ;
        RECT 8.915 229.570 9.295 236.730 ;
        RECT 24.375 229.570 24.755 236.730 ;
        RECT 47.675 234.335 49.950 234.845 ;
        RECT 52.575 234.335 54.875 234.845 ;
        RECT 57.170 234.335 59.450 234.845 ;
        RECT 86.295 234.355 88.570 234.865 ;
        RECT 91.195 234.355 93.495 234.865 ;
        RECT 95.790 234.355 98.070 234.865 ;
        RECT 122.550 229.590 122.930 236.750 ;
        RECT 8.495 217.680 80.885 217.820 ;
        RECT 8.495 216.920 137.210 217.680 ;
        RECT 8.865 209.760 9.245 216.920 ;
        RECT 24.325 209.760 24.705 216.920 ;
        RECT 80.855 216.780 137.210 216.920 ;
        RECT 47.625 214.525 49.900 215.035 ;
        RECT 52.525 214.525 54.825 215.035 ;
        RECT 57.120 214.525 59.400 215.035 ;
        RECT 86.295 214.385 88.570 214.895 ;
        RECT 91.195 214.385 93.495 214.895 ;
        RECT 95.790 214.385 98.070 214.895 ;
        RECT 122.550 209.620 122.930 216.780 ;
        RECT 8.465 198.015 80.855 198.025 ;
        RECT 8.465 197.125 137.210 198.015 ;
        RECT 8.835 189.965 9.215 197.125 ;
        RECT 24.295 189.965 24.675 197.125 ;
        RECT 80.855 197.115 137.210 197.125 ;
        RECT 47.595 194.730 49.870 195.240 ;
        RECT 52.495 194.730 54.795 195.240 ;
        RECT 57.090 194.730 59.370 195.240 ;
        RECT 86.295 194.720 88.570 195.230 ;
        RECT 91.195 194.720 93.495 195.230 ;
        RECT 95.790 194.720 98.070 195.230 ;
        RECT 122.550 189.955 122.930 197.115 ;
        RECT 8.615 178.175 81.005 178.230 ;
        RECT 8.615 177.330 137.250 178.175 ;
        RECT 8.985 170.170 9.365 177.330 ;
        RECT 24.445 170.170 24.825 177.330 ;
        RECT 80.895 177.275 137.250 177.330 ;
        RECT 47.745 174.935 50.020 175.445 ;
        RECT 52.645 174.935 54.945 175.445 ;
        RECT 57.240 174.935 59.520 175.445 ;
        RECT 86.335 174.880 88.610 175.390 ;
        RECT 91.235 174.880 93.535 175.390 ;
        RECT 95.830 174.880 98.110 175.390 ;
        RECT 122.590 170.115 122.970 177.275 ;
        RECT 8.570 158.450 80.960 158.540 ;
        RECT 8.570 157.640 137.050 158.450 ;
        RECT 8.940 150.480 9.320 157.640 ;
        RECT 24.400 150.480 24.780 157.640 ;
        RECT 80.695 157.550 137.050 157.640 ;
        RECT 47.700 155.245 49.975 155.755 ;
        RECT 52.600 155.245 54.900 155.755 ;
        RECT 57.195 155.245 59.475 155.755 ;
        RECT 86.135 155.155 88.410 155.665 ;
        RECT 91.035 155.155 93.335 155.665 ;
        RECT 95.630 155.155 97.910 155.665 ;
        RECT 122.390 150.390 122.770 157.550 ;
        RECT 8.760 138.805 81.150 138.830 ;
        RECT 8.760 137.930 137.205 138.805 ;
        RECT 9.130 130.770 9.510 137.930 ;
        RECT 24.590 130.770 24.970 137.930 ;
        RECT 80.850 137.905 137.205 137.930 ;
        RECT 47.890 135.535 50.165 136.045 ;
        RECT 52.790 135.535 55.090 136.045 ;
        RECT 57.385 135.535 59.665 136.045 ;
        RECT 86.290 135.510 88.565 136.020 ;
        RECT 91.190 135.510 93.490 136.020 ;
        RECT 95.785 135.510 98.065 136.020 ;
        RECT 122.545 130.745 122.925 137.905 ;
        RECT 80.850 118.990 137.205 119.010 ;
        RECT 8.565 118.110 137.205 118.990 ;
        RECT 8.565 118.090 80.955 118.110 ;
        RECT 8.935 110.930 9.315 118.090 ;
        RECT 24.395 110.930 24.775 118.090 ;
        RECT 47.695 115.695 49.970 116.205 ;
        RECT 52.595 115.695 54.895 116.205 ;
        RECT 57.190 115.695 59.470 116.205 ;
        RECT 86.290 115.715 88.565 116.225 ;
        RECT 91.190 115.715 93.490 116.225 ;
        RECT 95.785 115.715 98.065 116.225 ;
        RECT 122.545 110.950 122.925 118.110 ;
        RECT 8.435 99.255 80.825 99.280 ;
        RECT 8.435 98.380 137.125 99.255 ;
        RECT 8.805 91.220 9.185 98.380 ;
        RECT 24.265 91.220 24.645 98.380 ;
        RECT 80.770 98.355 137.125 98.380 ;
        RECT 47.565 95.985 49.840 96.495 ;
        RECT 52.465 95.985 54.765 96.495 ;
        RECT 57.060 95.985 59.340 96.495 ;
        RECT 86.210 95.960 88.485 96.470 ;
        RECT 91.110 95.960 93.410 96.470 ;
        RECT 95.705 95.960 97.985 96.470 ;
        RECT 122.465 91.195 122.845 98.355 ;
        RECT 80.875 79.520 137.230 79.540 ;
        RECT 8.565 78.640 137.230 79.520 ;
        RECT 8.565 78.620 80.955 78.640 ;
        RECT 8.935 71.460 9.315 78.620 ;
        RECT 24.395 71.460 24.775 78.620 ;
        RECT 47.695 76.225 49.970 76.735 ;
        RECT 52.595 76.225 54.895 76.735 ;
        RECT 57.190 76.225 59.470 76.735 ;
        RECT 86.315 76.245 88.590 76.755 ;
        RECT 91.215 76.245 93.515 76.755 ;
        RECT 95.810 76.245 98.090 76.755 ;
        RECT 122.570 71.480 122.950 78.640 ;
        RECT 8.515 59.570 80.905 59.710 ;
        RECT 8.515 58.810 137.230 59.570 ;
        RECT 8.885 51.650 9.265 58.810 ;
        RECT 24.345 51.650 24.725 58.810 ;
        RECT 80.875 58.670 137.230 58.810 ;
        RECT 47.645 56.415 49.920 56.925 ;
        RECT 52.545 56.415 54.845 56.925 ;
        RECT 57.140 56.415 59.420 56.925 ;
        RECT 86.315 56.275 88.590 56.785 ;
        RECT 91.215 56.275 93.515 56.785 ;
        RECT 95.810 56.275 98.090 56.785 ;
        RECT 122.570 51.510 122.950 58.670 ;
        RECT 8.485 39.905 80.875 39.915 ;
        RECT 8.485 39.015 137.230 39.905 ;
        RECT 8.855 31.855 9.235 39.015 ;
        RECT 24.315 31.855 24.695 39.015 ;
        RECT 80.875 39.005 137.230 39.015 ;
        RECT 47.615 36.620 49.890 37.130 ;
        RECT 52.515 36.620 54.815 37.130 ;
        RECT 57.110 36.620 59.390 37.130 ;
        RECT 86.315 36.610 88.590 37.120 ;
        RECT 91.215 36.610 93.515 37.120 ;
        RECT 95.810 36.610 98.090 37.120 ;
        RECT 122.570 31.845 122.950 39.005 ;
        RECT 79.670 19.270 94.700 20.170 ;
        RECT 93.950 12.110 94.330 19.270 ;
      LAYER Metal2 ;
        RECT 49.395 333.075 49.870 336.125 ;
        RECT 54.350 332.985 54.760 336.080 ;
        RECT 58.930 332.960 59.340 336.055 ;
        RECT 49.350 313.385 49.825 316.435 ;
        RECT 54.305 313.295 54.715 316.390 ;
        RECT 58.885 313.270 59.295 316.365 ;
        RECT 49.540 293.675 50.015 296.725 ;
        RECT 54.495 293.585 54.905 296.680 ;
        RECT 59.075 293.560 59.485 296.655 ;
        RECT 49.345 273.835 49.820 276.885 ;
        RECT 54.300 273.745 54.710 276.840 ;
        RECT 58.880 273.720 59.290 276.815 ;
        RECT 49.215 254.125 49.690 257.175 ;
        RECT 54.170 254.035 54.580 257.130 ;
        RECT 58.750 254.010 59.160 257.105 ;
        RECT 49.345 234.365 49.820 237.415 ;
        RECT 54.300 234.275 54.710 237.370 ;
        RECT 58.880 234.250 59.290 237.345 ;
        RECT 49.295 214.555 49.770 217.605 ;
        RECT 54.250 214.465 54.660 217.560 ;
        RECT 58.830 214.440 59.240 217.535 ;
        RECT 49.265 194.760 49.740 197.810 ;
        RECT 54.220 194.670 54.630 197.765 ;
        RECT 58.800 194.645 59.210 197.740 ;
        RECT 49.415 174.965 49.890 178.015 ;
        RECT 54.370 174.875 54.780 177.970 ;
        RECT 58.950 174.850 59.360 177.945 ;
        RECT 49.370 155.275 49.845 158.325 ;
        RECT 54.325 155.185 54.735 158.280 ;
        RECT 58.905 155.160 59.315 158.255 ;
        RECT 49.560 135.565 50.035 138.615 ;
        RECT 54.515 135.475 54.925 138.570 ;
        RECT 59.095 135.450 59.505 138.545 ;
        RECT 49.365 115.725 49.840 118.775 ;
        RECT 54.320 115.635 54.730 118.730 ;
        RECT 58.900 115.610 59.310 118.705 ;
        RECT 49.235 96.015 49.710 99.065 ;
        RECT 54.190 95.925 54.600 99.020 ;
        RECT 58.770 95.900 59.180 98.995 ;
        RECT 49.365 76.255 49.840 79.305 ;
        RECT 54.320 76.165 54.730 79.260 ;
        RECT 58.900 76.140 59.310 79.235 ;
        RECT 49.315 56.445 49.790 59.495 ;
        RECT 54.270 56.355 54.680 59.450 ;
        RECT 58.850 56.330 59.260 59.425 ;
        RECT 49.285 36.650 49.760 39.700 ;
        RECT 54.240 36.560 54.650 39.655 ;
        RECT 58.820 36.535 59.230 39.630 ;
        RECT 79.675 19.270 80.090 336.340 ;
        RECT 87.970 333.020 88.470 336.070 ;
        RECT 92.940 332.930 93.350 336.025 ;
        RECT 97.520 332.905 97.930 336.000 ;
        RECT 87.770 313.295 88.270 316.345 ;
        RECT 92.740 313.205 93.150 316.300 ;
        RECT 97.320 313.180 97.730 316.275 ;
        RECT 87.925 293.650 88.425 296.700 ;
        RECT 92.895 293.560 93.305 296.655 ;
        RECT 97.475 293.535 97.885 296.630 ;
        RECT 87.925 273.855 88.425 276.905 ;
        RECT 92.895 273.765 93.305 276.860 ;
        RECT 97.475 273.740 97.885 276.835 ;
        RECT 87.845 254.100 88.345 257.150 ;
        RECT 92.815 254.010 93.225 257.105 ;
        RECT 97.395 253.985 97.805 257.080 ;
        RECT 87.950 234.385 88.450 237.435 ;
        RECT 92.920 234.295 93.330 237.390 ;
        RECT 97.500 234.270 97.910 237.365 ;
        RECT 87.950 214.415 88.450 217.465 ;
        RECT 92.920 214.325 93.330 217.420 ;
        RECT 97.500 214.300 97.910 217.395 ;
        RECT 87.950 194.750 88.450 197.800 ;
        RECT 92.920 194.660 93.330 197.755 ;
        RECT 97.500 194.635 97.910 197.730 ;
        RECT 87.990 174.910 88.490 177.960 ;
        RECT 92.960 174.820 93.370 177.915 ;
        RECT 97.540 174.795 97.950 177.890 ;
        RECT 87.790 155.185 88.290 158.235 ;
        RECT 92.760 155.095 93.170 158.190 ;
        RECT 97.340 155.070 97.750 158.165 ;
        RECT 87.945 135.540 88.445 138.590 ;
        RECT 92.915 135.450 93.325 138.545 ;
        RECT 97.495 135.425 97.905 138.520 ;
        RECT 87.945 115.745 88.445 118.795 ;
        RECT 92.915 115.655 93.325 118.750 ;
        RECT 97.495 115.630 97.905 118.725 ;
        RECT 87.865 95.990 88.365 99.040 ;
        RECT 92.835 95.900 93.245 98.995 ;
        RECT 97.415 95.875 97.825 98.970 ;
        RECT 87.970 76.275 88.470 79.325 ;
        RECT 92.940 76.185 93.350 79.280 ;
        RECT 97.520 76.160 97.930 79.255 ;
        RECT 87.970 56.305 88.470 59.355 ;
        RECT 92.940 56.215 93.350 59.310 ;
        RECT 97.520 56.190 97.930 59.285 ;
        RECT 87.970 36.640 88.470 39.690 ;
        RECT 92.940 36.550 93.350 39.645 ;
        RECT 97.520 36.525 97.930 39.620 ;
      LAYER Metal3 ;
        RECT 14.100 22.065 80.105 22.555 ;
      LAYER Metal4 ;
        RECT 14.620 20.765 15.270 22.555 ;
        RECT 9.445 9.715 20.650 20.765 ;
    END
  END VDD
  OBS
      LAYER Metal1 ;
        RECT 41.065 334.400 78.615 334.455 ;
        RECT 41.065 334.170 106.635 334.400 ;
        RECT 77.860 334.115 106.635 334.170 ;
        RECT 108.305 334.095 115.010 334.395 ;
        RECT 44.770 333.260 45.970 333.640 ;
        RECT 64.295 333.360 65.530 333.740 ;
        RECT 81.165 333.205 82.620 333.585 ;
        RECT 104.860 333.305 106.140 333.685 ;
        RECT 65.710 333.005 66.090 333.040 ;
        RECT 44.210 332.900 44.590 332.940 ;
        RECT 44.140 332.595 46.975 332.900 ;
        RECT 62.955 332.695 66.090 333.005 ;
        RECT 104.300 332.950 104.680 332.985 ;
        RECT 82.800 332.845 83.180 332.885 ;
        RECT 65.710 332.660 66.090 332.695 ;
        RECT 44.210 332.560 44.590 332.595 ;
        RECT 82.730 332.540 85.565 332.845 ;
        RECT 101.545 332.640 104.680 332.950 ;
        RECT 123.810 332.925 130.550 333.225 ;
        RECT 104.300 332.605 104.680 332.640 ;
        RECT 82.800 332.505 83.180 332.540 ;
        RECT 14.540 330.985 14.920 331.365 ;
        RECT 21.440 330.975 21.820 331.355 ;
        RECT 30.000 330.985 30.380 331.365 ;
        RECT 36.900 330.975 37.280 331.355 ;
        RECT 44.770 330.960 48.030 331.340 ;
        RECT 48.770 330.960 52.030 331.340 ;
        RECT 58.270 330.960 61.530 331.340 ;
        RECT 62.270 330.960 65.530 331.340 ;
        RECT 81.325 330.905 82.620 331.285 ;
        RECT 87.360 330.905 90.620 331.285 ;
        RECT 91.360 330.905 92.545 331.285 ;
        RECT 94.810 330.905 96.120 331.285 ;
        RECT 96.860 330.905 100.120 331.285 ;
        RECT 104.860 330.905 105.875 331.285 ;
        RECT 108.940 331.150 112.355 331.570 ;
        RECT 115.400 330.970 115.780 331.350 ;
        RECT 124.400 331.130 127.855 331.570 ;
        RECT 130.860 330.970 131.240 331.350 ;
        RECT 11.865 330.560 13.605 330.850 ;
        RECT 18.365 330.480 20.975 330.905 ;
        RECT 27.325 330.560 29.065 330.850 ;
        RECT 33.825 330.480 36.420 330.855 ;
        RECT 44.210 330.260 44.590 330.640 ;
        RECT 48.210 330.260 48.590 330.640 ;
        RECT 52.210 330.595 52.590 330.640 ;
        RECT 57.710 330.595 58.090 330.640 ;
        RECT 52.160 330.280 58.095 330.595 ;
        RECT 52.210 330.260 52.590 330.280 ;
        RECT 57.710 330.260 58.090 330.280 ;
        RECT 61.710 330.260 62.090 330.640 ;
        RECT 65.710 330.260 66.090 330.640 ;
        RECT 82.800 330.205 83.180 330.585 ;
        RECT 86.800 330.205 87.180 330.585 ;
        RECT 90.800 330.540 91.180 330.585 ;
        RECT 96.300 330.540 96.680 330.585 ;
        RECT 90.750 330.225 96.685 330.540 ;
        RECT 90.800 330.205 91.180 330.225 ;
        RECT 96.300 330.205 96.680 330.225 ;
        RECT 100.300 330.205 100.680 330.585 ;
        RECT 104.300 330.205 104.680 330.585 ;
        RECT 113.800 330.455 115.000 330.745 ;
        RECT 120.720 330.520 121.100 330.900 ;
        RECT 129.260 330.455 130.460 330.745 ;
        RECT 136.180 330.520 136.560 330.900 ;
        RECT 74.890 329.580 95.665 329.955 ;
        RECT 45.435 329.045 72.745 329.385 ;
        RECT 20.550 328.040 23.655 328.315 ;
        RECT 36.010 328.040 39.760 328.315 ;
        RECT 73.920 328.225 105.885 328.615 ;
        RECT 41.065 327.915 59.735 327.925 ;
        RECT 41.065 327.870 71.085 327.915 ;
        RECT 41.065 327.860 98.325 327.870 ;
        RECT 41.065 327.605 107.330 327.860 ;
        RECT 70.765 327.550 107.330 327.605 ;
        RECT 40.535 326.880 76.445 326.935 ;
        RECT 40.535 326.665 107.730 326.880 ;
        RECT 75.985 326.610 107.730 326.665 ;
        RECT 111.950 326.490 118.340 326.780 ;
        RECT 127.410 326.490 133.800 326.780 ;
        RECT 13.220 325.965 23.875 326.300 ;
        RECT 28.680 325.965 39.185 326.300 ;
        RECT 64.155 326.100 74.705 326.435 ;
        RECT 44.750 325.460 48.050 325.840 ;
        RECT 48.750 325.460 52.050 325.840 ;
        RECT 58.250 325.460 61.550 325.840 ;
        RECT 62.250 325.460 65.550 325.840 ;
        RECT 81.335 325.405 82.640 325.785 ;
        RECT 87.340 325.405 90.640 325.785 ;
        RECT 91.340 325.405 92.700 325.785 ;
        RECT 94.675 325.405 96.140 325.785 ;
        RECT 96.840 325.405 100.140 325.785 ;
        RECT 104.840 325.405 106.020 325.785 ;
        RECT 44.210 325.115 44.590 325.150 ;
        RECT 13.190 324.645 14.970 324.935 ;
        RECT 20.565 324.615 21.875 324.935 ;
        RECT 28.650 324.645 30.430 324.935 ;
        RECT 36.025 324.615 37.335 324.935 ;
        RECT 43.945 324.805 46.955 325.115 ;
        RECT 44.210 324.770 44.590 324.805 ;
        RECT 48.210 324.770 49.300 325.150 ;
        RECT 52.210 325.145 52.590 325.150 ;
        RECT 49.730 324.780 52.595 325.145 ;
        RECT 57.710 325.125 58.090 325.150 ;
        RECT 57.695 324.805 59.840 325.125 ;
        RECT 52.210 324.770 52.590 324.780 ;
        RECT 57.710 324.770 58.090 324.805 ;
        RECT 60.755 324.770 62.090 325.150 ;
        RECT 65.710 325.130 66.090 325.150 ;
        RECT 63.245 324.810 66.155 325.130 ;
        RECT 82.800 325.060 83.180 325.095 ;
        RECT 65.710 324.770 66.090 324.810 ;
        RECT 82.535 324.750 85.545 325.060 ;
        RECT 82.800 324.715 83.180 324.750 ;
        RECT 86.800 324.715 87.890 325.095 ;
        RECT 90.800 325.090 91.180 325.095 ;
        RECT 88.320 324.725 91.185 325.090 ;
        RECT 96.300 325.070 96.680 325.095 ;
        RECT 96.285 324.750 98.430 325.070 ;
        RECT 90.800 324.715 91.180 324.725 ;
        RECT 96.300 324.715 96.680 324.750 ;
        RECT 99.345 324.715 100.680 325.095 ;
        RECT 104.300 325.075 104.680 325.095 ;
        RECT 101.835 324.755 104.745 325.075 ;
        RECT 104.300 324.715 104.680 324.755 ;
        RECT 108.930 324.575 109.310 324.955 ;
        RECT 114.590 324.680 115.780 324.965 ;
        RECT 124.390 324.575 124.770 324.955 ;
        RECT 130.050 324.680 131.240 324.965 ;
        RECT 11.920 324.030 12.300 324.410 ;
        RECT 18.375 324.060 18.755 324.440 ;
        RECT 27.380 324.030 27.760 324.410 ;
        RECT 33.835 324.060 34.215 324.440 ;
        RECT 113.810 324.015 114.190 324.395 ;
        RECT 117.930 323.850 121.110 324.170 ;
        RECT 129.270 324.015 129.650 324.395 ;
        RECT 133.390 323.850 136.570 324.170 ;
        RECT 44.750 323.460 46.035 323.840 ;
        RECT 64.065 323.460 65.550 323.840 ;
        RECT 81.150 323.405 82.640 323.785 ;
        RECT 104.840 323.405 105.915 323.785 ;
        RECT 44.210 322.770 45.300 323.150 ;
        RECT 48.695 322.775 61.545 323.110 ;
        RECT 65.710 323.105 66.090 323.150 ;
        RECT 64.975 322.805 66.285 323.105 ;
        RECT 65.710 322.770 66.090 322.805 ;
        RECT 82.800 322.715 83.890 323.095 ;
        RECT 87.285 322.720 100.135 323.055 ;
        RECT 104.300 323.050 104.680 323.095 ;
        RECT 103.565 322.750 104.875 323.050 ;
        RECT 123.670 322.765 127.820 323.035 ;
        RECT 104.300 322.715 104.680 322.750 ;
        RECT 41.065 322.220 74.145 322.260 ;
        RECT 41.065 321.910 106.310 322.220 ;
        RECT 73.360 321.855 106.310 321.910 ;
        RECT 108.105 321.845 112.365 322.200 ;
        RECT 41.020 314.675 78.570 314.765 ;
        RECT 41.020 314.480 106.435 314.675 ;
        RECT 77.660 314.390 106.435 314.480 ;
        RECT 108.105 314.370 114.810 314.670 ;
        RECT 44.725 313.570 45.925 313.950 ;
        RECT 64.250 313.670 65.485 314.050 ;
        RECT 80.965 313.480 82.420 313.860 ;
        RECT 104.660 313.580 105.940 313.960 ;
        RECT 65.665 313.315 66.045 313.350 ;
        RECT 44.165 313.210 44.545 313.250 ;
        RECT 44.095 312.905 46.930 313.210 ;
        RECT 62.910 313.005 66.045 313.315 ;
        RECT 104.100 313.225 104.480 313.260 ;
        RECT 82.600 313.120 82.980 313.160 ;
        RECT 65.665 312.970 66.045 313.005 ;
        RECT 44.165 312.870 44.545 312.905 ;
        RECT 82.530 312.815 85.365 313.120 ;
        RECT 101.345 312.915 104.480 313.225 ;
        RECT 123.610 313.200 130.350 313.500 ;
        RECT 104.100 312.880 104.480 312.915 ;
        RECT 82.600 312.780 82.980 312.815 ;
        RECT 14.495 311.295 14.875 311.675 ;
        RECT 21.395 311.285 21.775 311.665 ;
        RECT 26.210 311.495 29.615 311.935 ;
        RECT 29.955 311.295 30.335 311.675 ;
        RECT 32.670 311.335 33.050 311.715 ;
        RECT 36.855 311.285 37.235 311.665 ;
        RECT 44.725 311.270 47.985 311.650 ;
        RECT 48.725 311.270 51.985 311.650 ;
        RECT 58.225 311.270 61.485 311.650 ;
        RECT 62.225 311.270 65.485 311.650 ;
        RECT 11.820 310.870 13.560 311.160 ;
        RECT 18.320 310.790 20.930 311.215 ;
        RECT 27.280 310.870 29.020 311.160 ;
        RECT 31.070 310.820 32.270 311.110 ;
        RECT 33.780 310.790 36.375 311.165 ;
        RECT 37.990 310.885 38.370 311.265 ;
        RECT 81.125 311.180 82.420 311.560 ;
        RECT 87.160 311.180 90.420 311.560 ;
        RECT 91.160 311.180 92.345 311.560 ;
        RECT 94.610 311.180 95.920 311.560 ;
        RECT 96.660 311.180 99.920 311.560 ;
        RECT 104.660 311.180 105.675 311.560 ;
        RECT 108.740 311.425 112.155 311.845 ;
        RECT 112.485 311.205 112.865 311.585 ;
        RECT 115.200 311.245 115.580 311.625 ;
        RECT 119.385 311.195 119.765 311.575 ;
        RECT 124.200 311.405 127.655 311.845 ;
        RECT 130.660 311.245 131.040 311.625 ;
        RECT 44.165 310.570 44.545 310.950 ;
        RECT 48.165 310.570 48.545 310.950 ;
        RECT 52.165 310.905 52.545 310.950 ;
        RECT 57.665 310.905 58.045 310.950 ;
        RECT 52.115 310.590 58.050 310.905 ;
        RECT 52.165 310.570 52.545 310.590 ;
        RECT 57.665 310.570 58.045 310.590 ;
        RECT 61.665 310.570 62.045 310.950 ;
        RECT 65.665 310.570 66.045 310.950 ;
        RECT 82.600 310.480 82.980 310.860 ;
        RECT 86.600 310.480 86.980 310.860 ;
        RECT 90.600 310.815 90.980 310.860 ;
        RECT 96.100 310.815 96.480 310.860 ;
        RECT 90.550 310.500 96.485 310.815 ;
        RECT 90.600 310.480 90.980 310.500 ;
        RECT 96.100 310.480 96.480 310.500 ;
        RECT 100.100 310.480 100.480 310.860 ;
        RECT 104.100 310.480 104.480 310.860 ;
        RECT 109.810 310.780 111.550 311.070 ;
        RECT 113.600 310.730 114.800 311.020 ;
        RECT 116.310 310.690 118.940 311.145 ;
        RECT 120.520 310.795 120.900 311.175 ;
        RECT 129.060 310.730 130.260 311.020 ;
        RECT 135.980 310.795 136.360 311.175 ;
        RECT 74.690 309.855 95.465 310.230 ;
        RECT 123.015 310.020 138.935 310.320 ;
        RECT 45.390 309.355 72.700 309.695 ;
        RECT 123.550 309.275 140.495 309.575 ;
        RECT 25.005 308.650 32.265 308.950 ;
        RECT 20.505 308.350 23.610 308.625 ;
        RECT 25.560 308.115 29.645 308.385 ;
        RECT 35.965 308.350 39.715 308.625 ;
        RECT 73.720 308.500 105.685 308.890 ;
        RECT 118.495 308.260 121.625 308.535 ;
        RECT 41.020 308.225 59.690 308.235 ;
        RECT 41.020 308.145 71.040 308.225 ;
        RECT 41.020 308.135 98.125 308.145 ;
        RECT 41.020 307.915 107.130 308.135 ;
        RECT 70.565 307.825 107.130 307.915 ;
        RECT 124.745 307.365 128.875 307.665 ;
        RECT 131.250 307.315 135.750 307.625 ;
        RECT 40.490 307.155 76.400 307.245 ;
        RECT 29.220 306.855 35.610 307.145 ;
        RECT 40.490 306.975 107.530 307.155 ;
        RECT 75.785 306.885 107.530 306.975 ;
        RECT 111.750 306.765 118.140 307.055 ;
        RECT 127.210 306.765 133.600 307.055 ;
        RECT 13.175 306.275 23.830 306.610 ;
        RECT 28.635 306.275 39.140 306.610 ;
        RECT 64.110 306.410 74.660 306.745 ;
        RECT 111.165 306.185 121.645 306.520 ;
        RECT 44.705 305.770 48.005 306.150 ;
        RECT 48.705 305.770 52.005 306.150 ;
        RECT 58.205 305.770 61.505 306.150 ;
        RECT 62.205 305.770 65.505 306.150 ;
        RECT 81.135 305.680 82.440 306.060 ;
        RECT 87.140 305.680 90.440 306.060 ;
        RECT 91.140 305.680 92.500 306.060 ;
        RECT 94.475 305.680 95.940 306.060 ;
        RECT 96.640 305.680 99.940 306.060 ;
        RECT 104.640 305.680 105.820 306.060 ;
        RECT 125.975 305.600 128.895 305.900 ;
        RECT 132.440 305.585 135.810 305.885 ;
        RECT 44.165 305.425 44.545 305.460 ;
        RECT 13.145 304.955 14.925 305.245 ;
        RECT 20.520 304.925 21.830 305.245 ;
        RECT 26.200 304.940 26.580 305.320 ;
        RECT 28.605 304.955 30.385 305.245 ;
        RECT 31.860 305.045 33.050 305.330 ;
        RECT 35.980 304.925 37.290 305.245 ;
        RECT 43.900 305.115 46.910 305.425 ;
        RECT 44.165 305.080 44.545 305.115 ;
        RECT 48.165 305.080 49.255 305.460 ;
        RECT 52.165 305.455 52.545 305.460 ;
        RECT 49.685 305.090 52.550 305.455 ;
        RECT 57.665 305.435 58.045 305.460 ;
        RECT 57.650 305.115 59.795 305.435 ;
        RECT 52.165 305.080 52.545 305.090 ;
        RECT 57.665 305.080 58.045 305.115 ;
        RECT 60.710 305.080 62.045 305.460 ;
        RECT 65.665 305.440 66.045 305.460 ;
        RECT 63.200 305.120 66.110 305.440 ;
        RECT 82.600 305.335 82.980 305.370 ;
        RECT 65.665 305.080 66.045 305.120 ;
        RECT 82.335 305.025 85.345 305.335 ;
        RECT 82.600 304.990 82.980 305.025 ;
        RECT 86.600 304.990 87.690 305.370 ;
        RECT 90.600 305.365 90.980 305.370 ;
        RECT 88.120 305.000 90.985 305.365 ;
        RECT 96.100 305.345 96.480 305.370 ;
        RECT 96.085 305.025 98.230 305.345 ;
        RECT 90.600 304.990 90.980 305.000 ;
        RECT 96.100 304.990 96.480 305.025 ;
        RECT 99.145 304.990 100.480 305.370 ;
        RECT 104.100 305.350 104.480 305.370 ;
        RECT 101.635 305.030 104.545 305.350 ;
        RECT 104.100 304.990 104.480 305.030 ;
        RECT 108.730 304.850 109.110 305.230 ;
        RECT 111.135 304.865 112.915 305.155 ;
        RECT 114.390 304.955 115.580 305.240 ;
        RECT 118.510 304.835 119.820 305.155 ;
        RECT 124.190 304.850 124.570 305.230 ;
        RECT 129.850 304.955 131.040 305.240 ;
        RECT 11.875 304.340 12.255 304.720 ;
        RECT 18.330 304.370 18.710 304.750 ;
        RECT 27.335 304.340 27.715 304.720 ;
        RECT 31.080 304.380 31.460 304.760 ;
        RECT 33.790 304.370 34.170 304.750 ;
        RECT 35.200 304.215 38.380 304.535 ;
        RECT 109.865 304.250 110.245 304.630 ;
        RECT 113.610 304.290 113.990 304.670 ;
        RECT 116.320 304.280 116.700 304.660 ;
        RECT 44.705 303.770 45.990 304.150 ;
        RECT 64.020 303.770 65.505 304.150 ;
        RECT 117.730 304.125 120.910 304.445 ;
        RECT 129.070 304.290 129.450 304.670 ;
        RECT 133.190 304.125 136.370 304.445 ;
        RECT 80.950 303.680 82.440 304.060 ;
        RECT 104.640 303.680 105.715 304.060 ;
        RECT 44.165 303.080 45.255 303.460 ;
        RECT 48.650 303.085 61.500 303.420 ;
        RECT 65.665 303.415 66.045 303.460 ;
        RECT 64.930 303.115 66.240 303.415 ;
        RECT 65.665 303.080 66.045 303.115 ;
        RECT 82.600 302.990 83.690 303.370 ;
        RECT 87.085 302.995 99.935 303.330 ;
        RECT 104.100 303.325 104.480 303.370 ;
        RECT 103.365 303.025 104.675 303.325 ;
        RECT 123.470 303.040 127.620 303.310 ;
        RECT 104.100 302.990 104.480 303.025 ;
        RECT 41.020 302.495 74.100 302.570 ;
        RECT 41.020 302.220 106.110 302.495 ;
        RECT 73.160 302.130 106.110 302.220 ;
        RECT 107.905 302.120 112.165 302.475 ;
        RECT 41.210 295.030 78.760 295.055 ;
        RECT 41.210 294.770 106.590 295.030 ;
        RECT 77.815 294.745 106.590 294.770 ;
        RECT 108.260 294.725 114.965 295.025 ;
        RECT 44.915 293.860 46.115 294.240 ;
        RECT 64.440 293.960 65.675 294.340 ;
        RECT 81.120 293.835 82.575 294.215 ;
        RECT 104.815 293.935 106.095 294.315 ;
        RECT 65.855 293.605 66.235 293.640 ;
        RECT 44.355 293.500 44.735 293.540 ;
        RECT 44.285 293.195 47.120 293.500 ;
        RECT 63.100 293.295 66.235 293.605 ;
        RECT 104.255 293.580 104.635 293.615 ;
        RECT 82.755 293.475 83.135 293.515 ;
        RECT 65.855 293.260 66.235 293.295 ;
        RECT 44.355 293.160 44.735 293.195 ;
        RECT 82.685 293.170 85.520 293.475 ;
        RECT 101.500 293.270 104.635 293.580 ;
        RECT 123.765 293.555 130.505 293.855 ;
        RECT 104.255 293.235 104.635 293.270 ;
        RECT 82.755 293.135 83.135 293.170 ;
        RECT 14.685 291.585 15.065 291.965 ;
        RECT 21.585 291.575 21.965 291.955 ;
        RECT 26.400 291.785 29.805 292.225 ;
        RECT 30.145 291.585 30.525 291.965 ;
        RECT 32.860 291.625 33.240 292.005 ;
        RECT 37.045 291.575 37.425 291.955 ;
        RECT 44.915 291.560 48.175 291.940 ;
        RECT 48.915 291.560 52.175 291.940 ;
        RECT 58.415 291.560 61.675 291.940 ;
        RECT 62.415 291.560 65.675 291.940 ;
        RECT 12.010 291.160 13.750 291.450 ;
        RECT 18.510 291.080 21.120 291.505 ;
        RECT 27.470 291.160 29.210 291.450 ;
        RECT 31.260 291.110 32.460 291.400 ;
        RECT 33.970 291.080 36.565 291.455 ;
        RECT 38.180 291.175 38.560 291.555 ;
        RECT 81.280 291.535 82.575 291.915 ;
        RECT 87.315 291.535 90.575 291.915 ;
        RECT 91.315 291.535 92.500 291.915 ;
        RECT 94.765 291.535 96.075 291.915 ;
        RECT 96.815 291.535 100.075 291.915 ;
        RECT 104.815 291.535 105.830 291.915 ;
        RECT 108.895 291.780 112.310 292.200 ;
        RECT 112.640 291.560 113.020 291.940 ;
        RECT 115.355 291.600 115.735 291.980 ;
        RECT 119.540 291.550 119.920 291.930 ;
        RECT 124.355 291.760 127.810 292.200 ;
        RECT 130.815 291.600 131.195 291.980 ;
        RECT 44.355 290.860 44.735 291.240 ;
        RECT 48.355 290.860 48.735 291.240 ;
        RECT 52.355 291.195 52.735 291.240 ;
        RECT 57.855 291.195 58.235 291.240 ;
        RECT 52.305 290.880 58.240 291.195 ;
        RECT 52.355 290.860 52.735 290.880 ;
        RECT 57.855 290.860 58.235 290.880 ;
        RECT 61.855 290.860 62.235 291.240 ;
        RECT 65.855 290.860 66.235 291.240 ;
        RECT 82.755 290.835 83.135 291.215 ;
        RECT 86.755 290.835 87.135 291.215 ;
        RECT 90.755 291.170 91.135 291.215 ;
        RECT 96.255 291.170 96.635 291.215 ;
        RECT 90.705 290.855 96.640 291.170 ;
        RECT 90.755 290.835 91.135 290.855 ;
        RECT 96.255 290.835 96.635 290.855 ;
        RECT 100.255 290.835 100.635 291.215 ;
        RECT 104.255 290.835 104.635 291.215 ;
        RECT 109.965 291.135 111.705 291.425 ;
        RECT 113.755 291.085 114.955 291.375 ;
        RECT 116.465 291.045 119.095 291.500 ;
        RECT 120.675 291.150 121.055 291.530 ;
        RECT 129.215 291.085 130.415 291.375 ;
        RECT 136.135 291.150 136.515 291.530 ;
        RECT 74.845 290.210 95.620 290.585 ;
        RECT 123.170 290.375 139.090 290.675 ;
        RECT 45.580 289.645 72.890 289.985 ;
        RECT 123.705 289.630 140.650 289.930 ;
        RECT 25.195 288.940 32.455 289.240 ;
        RECT 20.695 288.640 23.800 288.915 ;
        RECT 25.750 288.405 29.835 288.675 ;
        RECT 36.155 288.640 39.905 288.915 ;
        RECT 73.875 288.855 105.840 289.245 ;
        RECT 118.650 288.615 121.780 288.890 ;
        RECT 41.210 288.515 59.880 288.525 ;
        RECT 41.210 288.500 71.230 288.515 ;
        RECT 41.210 288.490 98.280 288.500 ;
        RECT 41.210 288.205 107.285 288.490 ;
        RECT 70.720 288.180 107.285 288.205 ;
        RECT 124.900 287.720 129.030 288.020 ;
        RECT 131.405 287.670 135.905 287.980 ;
        RECT 40.680 287.510 76.590 287.535 ;
        RECT 29.410 287.145 35.800 287.435 ;
        RECT 40.680 287.265 107.685 287.510 ;
        RECT 75.940 287.240 107.685 287.265 ;
        RECT 111.905 287.120 118.295 287.410 ;
        RECT 127.365 287.120 133.755 287.410 ;
        RECT 13.365 286.565 24.020 286.900 ;
        RECT 28.825 286.565 39.330 286.900 ;
        RECT 64.300 286.700 74.850 287.035 ;
        RECT 111.320 286.540 121.800 286.875 ;
        RECT 44.895 286.060 48.195 286.440 ;
        RECT 48.895 286.060 52.195 286.440 ;
        RECT 58.395 286.060 61.695 286.440 ;
        RECT 62.395 286.060 65.695 286.440 ;
        RECT 81.290 286.035 82.595 286.415 ;
        RECT 87.295 286.035 90.595 286.415 ;
        RECT 91.295 286.035 92.655 286.415 ;
        RECT 94.630 286.035 96.095 286.415 ;
        RECT 96.795 286.035 100.095 286.415 ;
        RECT 104.795 286.035 105.975 286.415 ;
        RECT 126.130 285.955 129.050 286.255 ;
        RECT 132.595 285.940 135.965 286.240 ;
        RECT 44.355 285.715 44.735 285.750 ;
        RECT 13.335 285.245 15.115 285.535 ;
        RECT 20.710 285.215 22.020 285.535 ;
        RECT 26.390 285.230 26.770 285.610 ;
        RECT 28.795 285.245 30.575 285.535 ;
        RECT 32.050 285.335 33.240 285.620 ;
        RECT 36.170 285.215 37.480 285.535 ;
        RECT 44.090 285.405 47.100 285.715 ;
        RECT 44.355 285.370 44.735 285.405 ;
        RECT 48.355 285.370 49.445 285.750 ;
        RECT 52.355 285.745 52.735 285.750 ;
        RECT 49.875 285.380 52.740 285.745 ;
        RECT 57.855 285.725 58.235 285.750 ;
        RECT 57.840 285.405 59.985 285.725 ;
        RECT 52.355 285.370 52.735 285.380 ;
        RECT 57.855 285.370 58.235 285.405 ;
        RECT 60.900 285.370 62.235 285.750 ;
        RECT 65.855 285.730 66.235 285.750 ;
        RECT 63.390 285.410 66.300 285.730 ;
        RECT 82.755 285.690 83.135 285.725 ;
        RECT 65.855 285.370 66.235 285.410 ;
        RECT 82.490 285.380 85.500 285.690 ;
        RECT 82.755 285.345 83.135 285.380 ;
        RECT 86.755 285.345 87.845 285.725 ;
        RECT 90.755 285.720 91.135 285.725 ;
        RECT 88.275 285.355 91.140 285.720 ;
        RECT 96.255 285.700 96.635 285.725 ;
        RECT 96.240 285.380 98.385 285.700 ;
        RECT 90.755 285.345 91.135 285.355 ;
        RECT 96.255 285.345 96.635 285.380 ;
        RECT 99.300 285.345 100.635 285.725 ;
        RECT 104.255 285.705 104.635 285.725 ;
        RECT 101.790 285.385 104.700 285.705 ;
        RECT 104.255 285.345 104.635 285.385 ;
        RECT 108.885 285.205 109.265 285.585 ;
        RECT 111.290 285.220 113.070 285.510 ;
        RECT 114.545 285.310 115.735 285.595 ;
        RECT 118.665 285.190 119.975 285.510 ;
        RECT 124.345 285.205 124.725 285.585 ;
        RECT 130.005 285.310 131.195 285.595 ;
        RECT 12.065 284.630 12.445 285.010 ;
        RECT 18.520 284.660 18.900 285.040 ;
        RECT 27.525 284.630 27.905 285.010 ;
        RECT 31.270 284.670 31.650 285.050 ;
        RECT 33.980 284.660 34.360 285.040 ;
        RECT 35.390 284.505 38.570 284.825 ;
        RECT 110.020 284.605 110.400 284.985 ;
        RECT 113.765 284.645 114.145 285.025 ;
        RECT 116.475 284.635 116.855 285.015 ;
        RECT 117.885 284.480 121.065 284.800 ;
        RECT 129.225 284.645 129.605 285.025 ;
        RECT 133.345 284.480 136.525 284.800 ;
        RECT 44.895 284.060 46.180 284.440 ;
        RECT 64.210 284.060 65.695 284.440 ;
        RECT 81.105 284.035 82.595 284.415 ;
        RECT 104.795 284.035 105.870 284.415 ;
        RECT 44.355 283.370 45.445 283.750 ;
        RECT 48.840 283.375 61.690 283.710 ;
        RECT 65.855 283.705 66.235 283.750 ;
        RECT 65.120 283.405 66.430 283.705 ;
        RECT 65.855 283.370 66.235 283.405 ;
        RECT 82.755 283.345 83.845 283.725 ;
        RECT 87.240 283.350 100.090 283.685 ;
        RECT 104.255 283.680 104.635 283.725 ;
        RECT 103.520 283.380 104.830 283.680 ;
        RECT 123.625 283.395 127.775 283.665 ;
        RECT 104.255 283.345 104.635 283.380 ;
        RECT 41.210 282.850 74.290 282.860 ;
        RECT 41.210 282.510 106.265 282.850 ;
        RECT 73.315 282.485 106.265 282.510 ;
        RECT 108.060 282.475 112.320 282.830 ;
        RECT 77.815 275.215 106.590 275.235 ;
        RECT 41.015 274.950 106.590 275.215 ;
        RECT 41.015 274.930 78.565 274.950 ;
        RECT 108.260 274.930 114.965 275.230 ;
        RECT 44.720 274.020 45.920 274.400 ;
        RECT 64.245 274.120 65.480 274.500 ;
        RECT 81.120 274.040 82.575 274.420 ;
        RECT 104.815 274.140 106.095 274.520 ;
        RECT 65.660 273.765 66.040 273.800 ;
        RECT 104.255 273.785 104.635 273.820 ;
        RECT 44.160 273.660 44.540 273.700 ;
        RECT 44.090 273.355 46.925 273.660 ;
        RECT 62.905 273.455 66.040 273.765 ;
        RECT 82.755 273.680 83.135 273.720 ;
        RECT 65.660 273.420 66.040 273.455 ;
        RECT 82.685 273.375 85.520 273.680 ;
        RECT 101.500 273.475 104.635 273.785 ;
        RECT 123.765 273.760 130.505 274.060 ;
        RECT 104.255 273.440 104.635 273.475 ;
        RECT 44.160 273.320 44.540 273.355 ;
        RECT 82.755 273.340 83.135 273.375 ;
        RECT 14.490 271.745 14.870 272.125 ;
        RECT 21.390 271.735 21.770 272.115 ;
        RECT 26.205 271.945 29.610 272.385 ;
        RECT 29.950 271.745 30.330 272.125 ;
        RECT 32.665 271.785 33.045 272.165 ;
        RECT 36.850 271.735 37.230 272.115 ;
        RECT 44.720 271.720 47.980 272.100 ;
        RECT 48.720 271.720 51.980 272.100 ;
        RECT 58.220 271.720 61.480 272.100 ;
        RECT 62.220 271.720 65.480 272.100 ;
        RECT 81.280 271.740 82.575 272.120 ;
        RECT 87.315 271.740 90.575 272.120 ;
        RECT 91.315 271.740 92.500 272.120 ;
        RECT 94.765 271.740 96.075 272.120 ;
        RECT 96.815 271.740 100.075 272.120 ;
        RECT 104.815 271.740 105.830 272.120 ;
        RECT 108.895 271.985 112.310 272.405 ;
        RECT 112.640 271.765 113.020 272.145 ;
        RECT 115.355 271.805 115.735 272.185 ;
        RECT 119.540 271.755 119.920 272.135 ;
        RECT 124.355 271.965 127.810 272.405 ;
        RECT 130.815 271.805 131.195 272.185 ;
        RECT 11.815 271.320 13.555 271.610 ;
        RECT 18.315 271.240 20.925 271.665 ;
        RECT 27.275 271.320 29.015 271.610 ;
        RECT 31.065 271.270 32.265 271.560 ;
        RECT 33.775 271.240 36.370 271.615 ;
        RECT 37.985 271.335 38.365 271.715 ;
        RECT 44.160 271.020 44.540 271.400 ;
        RECT 48.160 271.020 48.540 271.400 ;
        RECT 52.160 271.355 52.540 271.400 ;
        RECT 57.660 271.355 58.040 271.400 ;
        RECT 52.110 271.040 58.045 271.355 ;
        RECT 52.160 271.020 52.540 271.040 ;
        RECT 57.660 271.020 58.040 271.040 ;
        RECT 61.660 271.020 62.040 271.400 ;
        RECT 65.660 271.020 66.040 271.400 ;
        RECT 82.755 271.040 83.135 271.420 ;
        RECT 86.755 271.040 87.135 271.420 ;
        RECT 90.755 271.375 91.135 271.420 ;
        RECT 96.255 271.375 96.635 271.420 ;
        RECT 90.705 271.060 96.640 271.375 ;
        RECT 90.755 271.040 91.135 271.060 ;
        RECT 96.255 271.040 96.635 271.060 ;
        RECT 100.255 271.040 100.635 271.420 ;
        RECT 104.255 271.040 104.635 271.420 ;
        RECT 109.965 271.340 111.705 271.630 ;
        RECT 113.755 271.290 114.955 271.580 ;
        RECT 116.465 271.250 119.095 271.705 ;
        RECT 120.675 271.355 121.055 271.735 ;
        RECT 129.215 271.290 130.415 271.580 ;
        RECT 136.135 271.355 136.515 271.735 ;
        RECT 74.845 270.415 95.620 270.790 ;
        RECT 123.170 270.580 139.090 270.880 ;
        RECT 45.385 269.805 72.695 270.145 ;
        RECT 123.705 269.835 140.650 270.135 ;
        RECT 25.000 269.100 32.260 269.400 ;
        RECT 20.500 268.800 23.605 269.075 ;
        RECT 25.555 268.565 29.640 268.835 ;
        RECT 35.960 268.800 39.710 269.075 ;
        RECT 73.875 269.060 105.840 269.450 ;
        RECT 118.650 268.820 121.780 269.095 ;
        RECT 70.720 268.695 98.280 268.705 ;
        RECT 41.015 268.675 59.685 268.685 ;
        RECT 70.720 268.675 107.285 268.695 ;
        RECT 41.015 268.385 107.285 268.675 ;
        RECT 41.015 268.365 71.035 268.385 ;
        RECT 124.900 267.925 129.030 268.225 ;
        RECT 131.405 267.875 135.905 268.185 ;
        RECT 75.940 267.695 107.685 267.715 ;
        RECT 29.215 267.305 35.605 267.595 ;
        RECT 40.485 267.445 107.685 267.695 ;
        RECT 40.485 267.425 76.395 267.445 ;
        RECT 111.905 267.325 118.295 267.615 ;
        RECT 127.365 267.325 133.755 267.615 ;
        RECT 13.170 266.725 23.825 267.060 ;
        RECT 28.630 266.725 39.135 267.060 ;
        RECT 64.105 266.860 74.655 267.195 ;
        RECT 111.320 266.745 121.800 267.080 ;
        RECT 44.700 266.220 48.000 266.600 ;
        RECT 48.700 266.220 52.000 266.600 ;
        RECT 58.200 266.220 61.500 266.600 ;
        RECT 62.200 266.220 65.500 266.600 ;
        RECT 81.290 266.240 82.595 266.620 ;
        RECT 87.295 266.240 90.595 266.620 ;
        RECT 91.295 266.240 92.655 266.620 ;
        RECT 94.630 266.240 96.095 266.620 ;
        RECT 96.795 266.240 100.095 266.620 ;
        RECT 104.795 266.240 105.975 266.620 ;
        RECT 126.130 266.160 129.050 266.460 ;
        RECT 132.595 266.145 135.965 266.445 ;
        RECT 44.160 265.875 44.540 265.910 ;
        RECT 13.140 265.405 14.920 265.695 ;
        RECT 20.515 265.375 21.825 265.695 ;
        RECT 26.195 265.390 26.575 265.770 ;
        RECT 28.600 265.405 30.380 265.695 ;
        RECT 31.855 265.495 33.045 265.780 ;
        RECT 35.975 265.375 37.285 265.695 ;
        RECT 43.895 265.565 46.905 265.875 ;
        RECT 44.160 265.530 44.540 265.565 ;
        RECT 48.160 265.530 49.250 265.910 ;
        RECT 52.160 265.905 52.540 265.910 ;
        RECT 49.680 265.540 52.545 265.905 ;
        RECT 57.660 265.885 58.040 265.910 ;
        RECT 57.645 265.565 59.790 265.885 ;
        RECT 52.160 265.530 52.540 265.540 ;
        RECT 57.660 265.530 58.040 265.565 ;
        RECT 60.705 265.530 62.040 265.910 ;
        RECT 65.660 265.890 66.040 265.910 ;
        RECT 82.755 265.895 83.135 265.930 ;
        RECT 63.195 265.570 66.105 265.890 ;
        RECT 82.490 265.585 85.500 265.895 ;
        RECT 65.660 265.530 66.040 265.570 ;
        RECT 82.755 265.550 83.135 265.585 ;
        RECT 86.755 265.550 87.845 265.930 ;
        RECT 90.755 265.925 91.135 265.930 ;
        RECT 88.275 265.560 91.140 265.925 ;
        RECT 96.255 265.905 96.635 265.930 ;
        RECT 96.240 265.585 98.385 265.905 ;
        RECT 90.755 265.550 91.135 265.560 ;
        RECT 96.255 265.550 96.635 265.585 ;
        RECT 99.300 265.550 100.635 265.930 ;
        RECT 104.255 265.910 104.635 265.930 ;
        RECT 101.790 265.590 104.700 265.910 ;
        RECT 104.255 265.550 104.635 265.590 ;
        RECT 108.885 265.410 109.265 265.790 ;
        RECT 111.290 265.425 113.070 265.715 ;
        RECT 114.545 265.515 115.735 265.800 ;
        RECT 118.665 265.395 119.975 265.715 ;
        RECT 124.345 265.410 124.725 265.790 ;
        RECT 130.005 265.515 131.195 265.800 ;
        RECT 11.870 264.790 12.250 265.170 ;
        RECT 18.325 264.820 18.705 265.200 ;
        RECT 27.330 264.790 27.710 265.170 ;
        RECT 31.075 264.830 31.455 265.210 ;
        RECT 33.785 264.820 34.165 265.200 ;
        RECT 35.195 264.665 38.375 264.985 ;
        RECT 110.020 264.810 110.400 265.190 ;
        RECT 113.765 264.850 114.145 265.230 ;
        RECT 116.475 264.840 116.855 265.220 ;
        RECT 117.885 264.685 121.065 265.005 ;
        RECT 129.225 264.850 129.605 265.230 ;
        RECT 133.345 264.685 136.525 265.005 ;
        RECT 44.700 264.220 45.985 264.600 ;
        RECT 64.015 264.220 65.500 264.600 ;
        RECT 81.105 264.240 82.595 264.620 ;
        RECT 104.795 264.240 105.870 264.620 ;
        RECT 44.160 263.530 45.250 263.910 ;
        RECT 48.645 263.535 61.495 263.870 ;
        RECT 65.660 263.865 66.040 263.910 ;
        RECT 64.925 263.565 66.235 263.865 ;
        RECT 65.660 263.530 66.040 263.565 ;
        RECT 82.755 263.550 83.845 263.930 ;
        RECT 87.240 263.555 100.090 263.890 ;
        RECT 104.255 263.885 104.635 263.930 ;
        RECT 103.520 263.585 104.830 263.885 ;
        RECT 123.625 263.600 127.775 263.870 ;
        RECT 104.255 263.550 104.635 263.585 ;
        RECT 73.315 263.020 106.265 263.055 ;
        RECT 41.015 262.690 106.265 263.020 ;
        RECT 41.015 262.670 74.095 262.690 ;
        RECT 108.060 262.680 112.320 263.035 ;
        RECT 40.885 255.480 78.435 255.505 ;
        RECT 40.885 255.220 106.510 255.480 ;
        RECT 77.735 255.195 106.510 255.220 ;
        RECT 108.180 255.175 114.885 255.475 ;
        RECT 44.590 254.310 45.790 254.690 ;
        RECT 64.115 254.410 65.350 254.790 ;
        RECT 81.040 254.285 82.495 254.665 ;
        RECT 104.735 254.385 106.015 254.765 ;
        RECT 65.530 254.055 65.910 254.090 ;
        RECT 44.030 253.950 44.410 253.990 ;
        RECT 43.960 253.645 46.795 253.950 ;
        RECT 62.775 253.745 65.910 254.055 ;
        RECT 104.175 254.030 104.555 254.065 ;
        RECT 82.675 253.925 83.055 253.965 ;
        RECT 65.530 253.710 65.910 253.745 ;
        RECT 44.030 253.610 44.410 253.645 ;
        RECT 82.605 253.620 85.440 253.925 ;
        RECT 101.420 253.720 104.555 254.030 ;
        RECT 123.685 254.005 130.425 254.305 ;
        RECT 104.175 253.685 104.555 253.720 ;
        RECT 82.675 253.585 83.055 253.620 ;
        RECT 14.360 252.035 14.740 252.415 ;
        RECT 21.260 252.025 21.640 252.405 ;
        RECT 26.075 252.235 29.480 252.675 ;
        RECT 29.820 252.035 30.200 252.415 ;
        RECT 32.535 252.075 32.915 252.455 ;
        RECT 36.720 252.025 37.100 252.405 ;
        RECT 44.590 252.010 47.850 252.390 ;
        RECT 48.590 252.010 51.850 252.390 ;
        RECT 58.090 252.010 61.350 252.390 ;
        RECT 62.090 252.010 65.350 252.390 ;
        RECT 11.685 251.610 13.425 251.900 ;
        RECT 18.185 251.530 20.795 251.955 ;
        RECT 27.145 251.610 28.885 251.900 ;
        RECT 30.935 251.560 32.135 251.850 ;
        RECT 33.645 251.530 36.240 251.905 ;
        RECT 37.855 251.625 38.235 252.005 ;
        RECT 81.200 251.985 82.495 252.365 ;
        RECT 87.235 251.985 90.495 252.365 ;
        RECT 91.235 251.985 92.420 252.365 ;
        RECT 94.685 251.985 95.995 252.365 ;
        RECT 96.735 251.985 99.995 252.365 ;
        RECT 104.735 251.985 105.750 252.365 ;
        RECT 108.815 252.230 112.230 252.650 ;
        RECT 112.560 252.010 112.940 252.390 ;
        RECT 115.275 252.050 115.655 252.430 ;
        RECT 119.460 252.000 119.840 252.380 ;
        RECT 124.275 252.210 127.730 252.650 ;
        RECT 130.735 252.050 131.115 252.430 ;
        RECT 44.030 251.310 44.410 251.690 ;
        RECT 48.030 251.310 48.410 251.690 ;
        RECT 52.030 251.645 52.410 251.690 ;
        RECT 57.530 251.645 57.910 251.690 ;
        RECT 51.980 251.330 57.915 251.645 ;
        RECT 52.030 251.310 52.410 251.330 ;
        RECT 57.530 251.310 57.910 251.330 ;
        RECT 61.530 251.310 61.910 251.690 ;
        RECT 65.530 251.310 65.910 251.690 ;
        RECT 82.675 251.285 83.055 251.665 ;
        RECT 86.675 251.285 87.055 251.665 ;
        RECT 90.675 251.620 91.055 251.665 ;
        RECT 96.175 251.620 96.555 251.665 ;
        RECT 90.625 251.305 96.560 251.620 ;
        RECT 90.675 251.285 91.055 251.305 ;
        RECT 96.175 251.285 96.555 251.305 ;
        RECT 100.175 251.285 100.555 251.665 ;
        RECT 104.175 251.285 104.555 251.665 ;
        RECT 109.885 251.585 111.625 251.875 ;
        RECT 113.675 251.535 114.875 251.825 ;
        RECT 116.385 251.495 119.015 251.950 ;
        RECT 120.595 251.600 120.975 251.980 ;
        RECT 129.135 251.535 130.335 251.825 ;
        RECT 136.055 251.600 136.435 251.980 ;
        RECT 74.765 250.660 95.540 251.035 ;
        RECT 123.090 250.825 139.010 251.125 ;
        RECT 45.255 250.095 72.565 250.435 ;
        RECT 123.625 250.080 140.570 250.380 ;
        RECT 24.870 249.390 32.130 249.690 ;
        RECT 20.370 249.090 23.475 249.365 ;
        RECT 25.425 248.855 29.510 249.125 ;
        RECT 35.830 249.090 39.580 249.365 ;
        RECT 73.795 249.305 105.760 249.695 ;
        RECT 118.570 249.065 121.700 249.340 ;
        RECT 40.885 248.965 59.555 248.975 ;
        RECT 40.885 248.950 70.905 248.965 ;
        RECT 40.885 248.940 98.200 248.950 ;
        RECT 40.885 248.655 107.205 248.940 ;
        RECT 70.640 248.630 107.205 248.655 ;
        RECT 124.820 248.170 128.950 248.470 ;
        RECT 131.325 248.120 135.825 248.430 ;
        RECT 40.355 247.960 76.265 247.985 ;
        RECT 29.085 247.595 35.475 247.885 ;
        RECT 40.355 247.715 107.605 247.960 ;
        RECT 75.860 247.690 107.605 247.715 ;
        RECT 111.825 247.570 118.215 247.860 ;
        RECT 127.285 247.570 133.675 247.860 ;
        RECT 13.040 247.015 23.695 247.350 ;
        RECT 28.500 247.015 39.005 247.350 ;
        RECT 63.975 247.150 74.525 247.485 ;
        RECT 111.240 246.990 121.720 247.325 ;
        RECT 44.570 246.510 47.870 246.890 ;
        RECT 48.570 246.510 51.870 246.890 ;
        RECT 58.070 246.510 61.370 246.890 ;
        RECT 62.070 246.510 65.370 246.890 ;
        RECT 81.210 246.485 82.515 246.865 ;
        RECT 87.215 246.485 90.515 246.865 ;
        RECT 91.215 246.485 92.575 246.865 ;
        RECT 94.550 246.485 96.015 246.865 ;
        RECT 96.715 246.485 100.015 246.865 ;
        RECT 104.715 246.485 105.895 246.865 ;
        RECT 126.050 246.405 128.970 246.705 ;
        RECT 132.515 246.390 135.885 246.690 ;
        RECT 44.030 246.165 44.410 246.200 ;
        RECT 13.010 245.695 14.790 245.985 ;
        RECT 20.385 245.665 21.695 245.985 ;
        RECT 26.065 245.680 26.445 246.060 ;
        RECT 28.470 245.695 30.250 245.985 ;
        RECT 31.725 245.785 32.915 246.070 ;
        RECT 35.845 245.665 37.155 245.985 ;
        RECT 43.765 245.855 46.775 246.165 ;
        RECT 44.030 245.820 44.410 245.855 ;
        RECT 48.030 245.820 49.120 246.200 ;
        RECT 52.030 246.195 52.410 246.200 ;
        RECT 49.550 245.830 52.415 246.195 ;
        RECT 57.530 246.175 57.910 246.200 ;
        RECT 57.515 245.855 59.660 246.175 ;
        RECT 52.030 245.820 52.410 245.830 ;
        RECT 57.530 245.820 57.910 245.855 ;
        RECT 60.575 245.820 61.910 246.200 ;
        RECT 65.530 246.180 65.910 246.200 ;
        RECT 63.065 245.860 65.975 246.180 ;
        RECT 82.675 246.140 83.055 246.175 ;
        RECT 65.530 245.820 65.910 245.860 ;
        RECT 82.410 245.830 85.420 246.140 ;
        RECT 82.675 245.795 83.055 245.830 ;
        RECT 86.675 245.795 87.765 246.175 ;
        RECT 90.675 246.170 91.055 246.175 ;
        RECT 88.195 245.805 91.060 246.170 ;
        RECT 96.175 246.150 96.555 246.175 ;
        RECT 96.160 245.830 98.305 246.150 ;
        RECT 90.675 245.795 91.055 245.805 ;
        RECT 96.175 245.795 96.555 245.830 ;
        RECT 99.220 245.795 100.555 246.175 ;
        RECT 104.175 246.155 104.555 246.175 ;
        RECT 101.710 245.835 104.620 246.155 ;
        RECT 104.175 245.795 104.555 245.835 ;
        RECT 108.805 245.655 109.185 246.035 ;
        RECT 111.210 245.670 112.990 245.960 ;
        RECT 114.465 245.760 115.655 246.045 ;
        RECT 118.585 245.640 119.895 245.960 ;
        RECT 124.265 245.655 124.645 246.035 ;
        RECT 129.925 245.760 131.115 246.045 ;
        RECT 11.740 245.080 12.120 245.460 ;
        RECT 18.195 245.110 18.575 245.490 ;
        RECT 27.200 245.080 27.580 245.460 ;
        RECT 30.945 245.120 31.325 245.500 ;
        RECT 33.655 245.110 34.035 245.490 ;
        RECT 35.065 244.955 38.245 245.275 ;
        RECT 109.940 245.055 110.320 245.435 ;
        RECT 113.685 245.095 114.065 245.475 ;
        RECT 116.395 245.085 116.775 245.465 ;
        RECT 117.805 244.930 120.985 245.250 ;
        RECT 129.145 245.095 129.525 245.475 ;
        RECT 133.265 244.930 136.445 245.250 ;
        RECT 44.570 244.510 45.855 244.890 ;
        RECT 63.885 244.510 65.370 244.890 ;
        RECT 81.025 244.485 82.515 244.865 ;
        RECT 104.715 244.485 105.790 244.865 ;
        RECT 44.030 243.820 45.120 244.200 ;
        RECT 48.515 243.825 61.365 244.160 ;
        RECT 65.530 244.155 65.910 244.200 ;
        RECT 64.795 243.855 66.105 244.155 ;
        RECT 65.530 243.820 65.910 243.855 ;
        RECT 82.675 243.795 83.765 244.175 ;
        RECT 87.160 243.800 100.010 244.135 ;
        RECT 104.175 244.130 104.555 244.175 ;
        RECT 103.440 243.830 104.750 244.130 ;
        RECT 123.545 243.845 127.695 244.115 ;
        RECT 104.175 243.795 104.555 243.830 ;
        RECT 40.885 243.300 73.965 243.310 ;
        RECT 40.885 242.960 106.185 243.300 ;
        RECT 73.235 242.935 106.185 242.960 ;
        RECT 107.980 242.925 112.240 243.280 ;
        RECT 77.840 235.745 106.615 235.765 ;
        RECT 41.015 235.480 106.615 235.745 ;
        RECT 41.015 235.460 78.565 235.480 ;
        RECT 108.285 235.460 114.990 235.760 ;
        RECT 44.720 234.550 45.920 234.930 ;
        RECT 64.245 234.650 65.480 235.030 ;
        RECT 81.145 234.570 82.600 234.950 ;
        RECT 104.840 234.670 106.120 235.050 ;
        RECT 65.660 234.295 66.040 234.330 ;
        RECT 104.280 234.315 104.660 234.350 ;
        RECT 44.160 234.190 44.540 234.230 ;
        RECT 44.090 233.885 46.925 234.190 ;
        RECT 62.905 233.985 66.040 234.295 ;
        RECT 82.780 234.210 83.160 234.250 ;
        RECT 65.660 233.950 66.040 233.985 ;
        RECT 82.710 233.905 85.545 234.210 ;
        RECT 101.525 234.005 104.660 234.315 ;
        RECT 123.790 234.290 130.530 234.590 ;
        RECT 104.280 233.970 104.660 234.005 ;
        RECT 44.160 233.850 44.540 233.885 ;
        RECT 82.780 233.870 83.160 233.905 ;
        RECT 14.490 232.275 14.870 232.655 ;
        RECT 21.390 232.265 21.770 232.645 ;
        RECT 26.205 232.475 29.610 232.915 ;
        RECT 29.950 232.275 30.330 232.655 ;
        RECT 32.665 232.315 33.045 232.695 ;
        RECT 36.850 232.265 37.230 232.645 ;
        RECT 44.720 232.250 47.980 232.630 ;
        RECT 48.720 232.250 51.980 232.630 ;
        RECT 58.220 232.250 61.480 232.630 ;
        RECT 62.220 232.250 65.480 232.630 ;
        RECT 81.305 232.270 82.600 232.650 ;
        RECT 87.340 232.270 90.600 232.650 ;
        RECT 91.340 232.270 92.525 232.650 ;
        RECT 94.790 232.270 96.100 232.650 ;
        RECT 96.840 232.270 100.100 232.650 ;
        RECT 104.840 232.270 105.855 232.650 ;
        RECT 108.920 232.515 112.335 232.935 ;
        RECT 112.665 232.295 113.045 232.675 ;
        RECT 115.380 232.335 115.760 232.715 ;
        RECT 119.565 232.285 119.945 232.665 ;
        RECT 124.380 232.495 127.835 232.935 ;
        RECT 130.840 232.335 131.220 232.715 ;
        RECT 11.815 231.850 13.555 232.140 ;
        RECT 18.315 231.770 20.925 232.195 ;
        RECT 27.275 231.850 29.015 232.140 ;
        RECT 31.065 231.800 32.265 232.090 ;
        RECT 33.775 231.770 36.370 232.145 ;
        RECT 37.985 231.865 38.365 232.245 ;
        RECT 44.160 231.550 44.540 231.930 ;
        RECT 48.160 231.550 48.540 231.930 ;
        RECT 52.160 231.885 52.540 231.930 ;
        RECT 57.660 231.885 58.040 231.930 ;
        RECT 52.110 231.570 58.045 231.885 ;
        RECT 52.160 231.550 52.540 231.570 ;
        RECT 57.660 231.550 58.040 231.570 ;
        RECT 61.660 231.550 62.040 231.930 ;
        RECT 65.660 231.550 66.040 231.930 ;
        RECT 82.780 231.570 83.160 231.950 ;
        RECT 86.780 231.570 87.160 231.950 ;
        RECT 90.780 231.905 91.160 231.950 ;
        RECT 96.280 231.905 96.660 231.950 ;
        RECT 90.730 231.590 96.665 231.905 ;
        RECT 90.780 231.570 91.160 231.590 ;
        RECT 96.280 231.570 96.660 231.590 ;
        RECT 100.280 231.570 100.660 231.950 ;
        RECT 104.280 231.570 104.660 231.950 ;
        RECT 109.990 231.870 111.730 232.160 ;
        RECT 113.780 231.820 114.980 232.110 ;
        RECT 116.490 231.780 119.120 232.235 ;
        RECT 120.700 231.885 121.080 232.265 ;
        RECT 129.240 231.820 130.440 232.110 ;
        RECT 136.160 231.885 136.540 232.265 ;
        RECT 74.870 230.945 95.645 231.320 ;
        RECT 123.195 231.110 139.115 231.410 ;
        RECT 45.385 230.335 72.695 230.675 ;
        RECT 123.730 230.365 140.675 230.665 ;
        RECT 25.000 229.630 32.260 229.930 ;
        RECT 20.500 229.330 23.605 229.605 ;
        RECT 25.555 229.095 29.640 229.365 ;
        RECT 35.960 229.330 39.710 229.605 ;
        RECT 73.900 229.590 105.865 229.980 ;
        RECT 118.675 229.350 121.805 229.625 ;
        RECT 70.745 229.225 98.305 229.235 ;
        RECT 41.015 229.205 59.685 229.215 ;
        RECT 70.745 229.205 107.310 229.225 ;
        RECT 41.015 228.915 107.310 229.205 ;
        RECT 41.015 228.895 71.035 228.915 ;
        RECT 124.925 228.455 129.055 228.755 ;
        RECT 131.430 228.405 135.930 228.715 ;
        RECT 75.965 228.225 107.710 228.245 ;
        RECT 29.215 227.835 35.605 228.125 ;
        RECT 40.485 227.975 107.710 228.225 ;
        RECT 40.485 227.955 76.395 227.975 ;
        RECT 111.930 227.855 118.320 228.145 ;
        RECT 127.390 227.855 133.780 228.145 ;
        RECT 13.170 227.255 23.825 227.590 ;
        RECT 28.630 227.255 39.135 227.590 ;
        RECT 64.105 227.390 74.655 227.725 ;
        RECT 111.345 227.275 121.825 227.610 ;
        RECT 44.700 226.750 48.000 227.130 ;
        RECT 48.700 226.750 52.000 227.130 ;
        RECT 58.200 226.750 61.500 227.130 ;
        RECT 62.200 226.750 65.500 227.130 ;
        RECT 81.315 226.770 82.620 227.150 ;
        RECT 87.320 226.770 90.620 227.150 ;
        RECT 91.320 226.770 92.680 227.150 ;
        RECT 94.655 226.770 96.120 227.150 ;
        RECT 96.820 226.770 100.120 227.150 ;
        RECT 104.820 226.770 106.000 227.150 ;
        RECT 126.155 226.690 129.075 226.990 ;
        RECT 132.620 226.675 135.990 226.975 ;
        RECT 44.160 226.405 44.540 226.440 ;
        RECT 13.140 225.935 14.920 226.225 ;
        RECT 20.515 225.905 21.825 226.225 ;
        RECT 26.195 225.920 26.575 226.300 ;
        RECT 28.600 225.935 30.380 226.225 ;
        RECT 31.855 226.025 33.045 226.310 ;
        RECT 35.975 225.905 37.285 226.225 ;
        RECT 43.895 226.095 46.905 226.405 ;
        RECT 44.160 226.060 44.540 226.095 ;
        RECT 48.160 226.060 49.250 226.440 ;
        RECT 52.160 226.435 52.540 226.440 ;
        RECT 49.680 226.070 52.545 226.435 ;
        RECT 57.660 226.415 58.040 226.440 ;
        RECT 57.645 226.095 59.790 226.415 ;
        RECT 52.160 226.060 52.540 226.070 ;
        RECT 57.660 226.060 58.040 226.095 ;
        RECT 60.705 226.060 62.040 226.440 ;
        RECT 65.660 226.420 66.040 226.440 ;
        RECT 82.780 226.425 83.160 226.460 ;
        RECT 63.195 226.100 66.105 226.420 ;
        RECT 82.515 226.115 85.525 226.425 ;
        RECT 65.660 226.060 66.040 226.100 ;
        RECT 82.780 226.080 83.160 226.115 ;
        RECT 86.780 226.080 87.870 226.460 ;
        RECT 90.780 226.455 91.160 226.460 ;
        RECT 88.300 226.090 91.165 226.455 ;
        RECT 96.280 226.435 96.660 226.460 ;
        RECT 96.265 226.115 98.410 226.435 ;
        RECT 90.780 226.080 91.160 226.090 ;
        RECT 96.280 226.080 96.660 226.115 ;
        RECT 99.325 226.080 100.660 226.460 ;
        RECT 104.280 226.440 104.660 226.460 ;
        RECT 101.815 226.120 104.725 226.440 ;
        RECT 104.280 226.080 104.660 226.120 ;
        RECT 108.910 225.940 109.290 226.320 ;
        RECT 111.315 225.955 113.095 226.245 ;
        RECT 114.570 226.045 115.760 226.330 ;
        RECT 118.690 225.925 120.000 226.245 ;
        RECT 124.370 225.940 124.750 226.320 ;
        RECT 130.030 226.045 131.220 226.330 ;
        RECT 11.870 225.320 12.250 225.700 ;
        RECT 18.325 225.350 18.705 225.730 ;
        RECT 27.330 225.320 27.710 225.700 ;
        RECT 31.075 225.360 31.455 225.740 ;
        RECT 33.785 225.350 34.165 225.730 ;
        RECT 35.195 225.195 38.375 225.515 ;
        RECT 110.045 225.340 110.425 225.720 ;
        RECT 113.790 225.380 114.170 225.760 ;
        RECT 116.500 225.370 116.880 225.750 ;
        RECT 117.910 225.215 121.090 225.535 ;
        RECT 129.250 225.380 129.630 225.760 ;
        RECT 133.370 225.215 136.550 225.535 ;
        RECT 44.700 224.750 45.985 225.130 ;
        RECT 64.015 224.750 65.500 225.130 ;
        RECT 81.130 224.770 82.620 225.150 ;
        RECT 104.820 224.770 105.895 225.150 ;
        RECT 44.160 224.060 45.250 224.440 ;
        RECT 48.645 224.065 61.495 224.400 ;
        RECT 65.660 224.395 66.040 224.440 ;
        RECT 64.925 224.095 66.235 224.395 ;
        RECT 65.660 224.060 66.040 224.095 ;
        RECT 82.780 224.080 83.870 224.460 ;
        RECT 87.265 224.085 100.115 224.420 ;
        RECT 104.280 224.415 104.660 224.460 ;
        RECT 103.545 224.115 104.855 224.415 ;
        RECT 123.650 224.130 127.800 224.400 ;
        RECT 104.280 224.080 104.660 224.115 ;
        RECT 73.340 223.550 106.290 223.585 ;
        RECT 41.015 223.220 106.290 223.550 ;
        RECT 41.015 223.200 74.095 223.220 ;
        RECT 108.085 223.210 112.345 223.565 ;
        RECT 40.965 215.795 78.515 215.935 ;
        RECT 40.965 215.650 106.615 215.795 ;
        RECT 77.840 215.510 106.615 215.650 ;
        RECT 108.285 215.490 114.990 215.790 ;
        RECT 44.670 214.740 45.870 215.120 ;
        RECT 64.195 214.840 65.430 215.220 ;
        RECT 81.145 214.600 82.600 214.980 ;
        RECT 104.840 214.700 106.120 215.080 ;
        RECT 65.610 214.485 65.990 214.520 ;
        RECT 44.110 214.380 44.490 214.420 ;
        RECT 44.040 214.075 46.875 214.380 ;
        RECT 62.855 214.175 65.990 214.485 ;
        RECT 104.280 214.345 104.660 214.380 ;
        RECT 82.780 214.240 83.160 214.280 ;
        RECT 65.610 214.140 65.990 214.175 ;
        RECT 44.110 214.040 44.490 214.075 ;
        RECT 82.710 213.935 85.545 214.240 ;
        RECT 101.525 214.035 104.660 214.345 ;
        RECT 123.790 214.320 130.530 214.620 ;
        RECT 104.280 214.000 104.660 214.035 ;
        RECT 82.780 213.900 83.160 213.935 ;
        RECT 14.440 212.465 14.820 212.845 ;
        RECT 21.340 212.455 21.720 212.835 ;
        RECT 26.155 212.665 29.560 213.105 ;
        RECT 29.900 212.465 30.280 212.845 ;
        RECT 32.615 212.505 32.995 212.885 ;
        RECT 36.800 212.455 37.180 212.835 ;
        RECT 44.670 212.440 47.930 212.820 ;
        RECT 48.670 212.440 51.930 212.820 ;
        RECT 58.170 212.440 61.430 212.820 ;
        RECT 62.170 212.440 65.430 212.820 ;
        RECT 11.765 212.040 13.505 212.330 ;
        RECT 18.265 211.960 20.875 212.385 ;
        RECT 27.225 212.040 28.965 212.330 ;
        RECT 31.015 211.990 32.215 212.280 ;
        RECT 33.725 211.960 36.320 212.335 ;
        RECT 37.935 212.055 38.315 212.435 ;
        RECT 81.305 212.300 82.600 212.680 ;
        RECT 87.340 212.300 90.600 212.680 ;
        RECT 91.340 212.300 92.525 212.680 ;
        RECT 94.790 212.300 96.100 212.680 ;
        RECT 96.840 212.300 100.100 212.680 ;
        RECT 104.840 212.300 105.855 212.680 ;
        RECT 108.920 212.545 112.335 212.965 ;
        RECT 112.665 212.325 113.045 212.705 ;
        RECT 115.380 212.365 115.760 212.745 ;
        RECT 119.565 212.315 119.945 212.695 ;
        RECT 124.380 212.525 127.835 212.965 ;
        RECT 130.840 212.365 131.220 212.745 ;
        RECT 44.110 211.740 44.490 212.120 ;
        RECT 48.110 211.740 48.490 212.120 ;
        RECT 52.110 212.075 52.490 212.120 ;
        RECT 57.610 212.075 57.990 212.120 ;
        RECT 52.060 211.760 57.995 212.075 ;
        RECT 52.110 211.740 52.490 211.760 ;
        RECT 57.610 211.740 57.990 211.760 ;
        RECT 61.610 211.740 61.990 212.120 ;
        RECT 65.610 211.740 65.990 212.120 ;
        RECT 82.780 211.600 83.160 211.980 ;
        RECT 86.780 211.600 87.160 211.980 ;
        RECT 90.780 211.935 91.160 211.980 ;
        RECT 96.280 211.935 96.660 211.980 ;
        RECT 90.730 211.620 96.665 211.935 ;
        RECT 90.780 211.600 91.160 211.620 ;
        RECT 96.280 211.600 96.660 211.620 ;
        RECT 100.280 211.600 100.660 211.980 ;
        RECT 104.280 211.600 104.660 211.980 ;
        RECT 109.990 211.900 111.730 212.190 ;
        RECT 113.780 211.850 114.980 212.140 ;
        RECT 116.490 211.810 119.120 212.265 ;
        RECT 120.700 211.915 121.080 212.295 ;
        RECT 129.240 211.850 130.440 212.140 ;
        RECT 136.160 211.915 136.540 212.295 ;
        RECT 74.870 210.975 95.645 211.350 ;
        RECT 123.195 211.140 139.115 211.440 ;
        RECT 45.335 210.525 72.645 210.865 ;
        RECT 123.730 210.395 140.675 210.695 ;
        RECT 24.950 209.820 32.210 210.120 ;
        RECT 20.450 209.520 23.555 209.795 ;
        RECT 25.505 209.285 29.590 209.555 ;
        RECT 35.910 209.520 39.660 209.795 ;
        RECT 73.900 209.620 105.865 210.010 ;
        RECT 40.965 209.395 59.635 209.405 ;
        RECT 40.965 209.265 70.985 209.395 ;
        RECT 118.675 209.380 121.805 209.655 ;
        RECT 40.965 209.255 98.305 209.265 ;
        RECT 40.965 209.085 107.310 209.255 ;
        RECT 70.745 208.945 107.310 209.085 ;
        RECT 124.925 208.485 129.055 208.785 ;
        RECT 131.430 208.435 135.930 208.745 ;
        RECT 29.165 208.025 35.555 208.315 ;
        RECT 40.435 208.275 76.345 208.415 ;
        RECT 40.435 208.145 107.710 208.275 ;
        RECT 75.965 208.005 107.710 208.145 ;
        RECT 13.120 207.445 23.775 207.780 ;
        RECT 28.580 207.445 39.085 207.780 ;
        RECT 64.055 207.580 74.605 207.915 ;
        RECT 111.930 207.885 118.320 208.175 ;
        RECT 127.390 207.885 133.780 208.175 ;
        RECT 44.650 206.940 47.950 207.320 ;
        RECT 48.650 206.940 51.950 207.320 ;
        RECT 58.150 206.940 61.450 207.320 ;
        RECT 62.150 206.940 65.450 207.320 ;
        RECT 111.345 207.305 121.825 207.640 ;
        RECT 81.315 206.800 82.620 207.180 ;
        RECT 87.320 206.800 90.620 207.180 ;
        RECT 91.320 206.800 92.680 207.180 ;
        RECT 94.655 206.800 96.120 207.180 ;
        RECT 96.820 206.800 100.120 207.180 ;
        RECT 104.820 206.800 106.000 207.180 ;
        RECT 126.155 206.720 129.075 207.020 ;
        RECT 132.620 206.705 135.990 207.005 ;
        RECT 44.110 206.595 44.490 206.630 ;
        RECT 13.090 206.125 14.870 206.415 ;
        RECT 20.465 206.095 21.775 206.415 ;
        RECT 26.145 206.110 26.525 206.490 ;
        RECT 28.550 206.125 30.330 206.415 ;
        RECT 31.805 206.215 32.995 206.500 ;
        RECT 35.925 206.095 37.235 206.415 ;
        RECT 43.845 206.285 46.855 206.595 ;
        RECT 44.110 206.250 44.490 206.285 ;
        RECT 48.110 206.250 49.200 206.630 ;
        RECT 52.110 206.625 52.490 206.630 ;
        RECT 49.630 206.260 52.495 206.625 ;
        RECT 57.610 206.605 57.990 206.630 ;
        RECT 57.595 206.285 59.740 206.605 ;
        RECT 52.110 206.250 52.490 206.260 ;
        RECT 57.610 206.250 57.990 206.285 ;
        RECT 60.655 206.250 61.990 206.630 ;
        RECT 65.610 206.610 65.990 206.630 ;
        RECT 63.145 206.290 66.055 206.610 ;
        RECT 82.780 206.455 83.160 206.490 ;
        RECT 65.610 206.250 65.990 206.290 ;
        RECT 82.515 206.145 85.525 206.455 ;
        RECT 82.780 206.110 83.160 206.145 ;
        RECT 86.780 206.110 87.870 206.490 ;
        RECT 90.780 206.485 91.160 206.490 ;
        RECT 88.300 206.120 91.165 206.485 ;
        RECT 96.280 206.465 96.660 206.490 ;
        RECT 96.265 206.145 98.410 206.465 ;
        RECT 90.780 206.110 91.160 206.120 ;
        RECT 96.280 206.110 96.660 206.145 ;
        RECT 99.325 206.110 100.660 206.490 ;
        RECT 104.280 206.470 104.660 206.490 ;
        RECT 101.815 206.150 104.725 206.470 ;
        RECT 104.280 206.110 104.660 206.150 ;
        RECT 108.910 205.970 109.290 206.350 ;
        RECT 111.315 205.985 113.095 206.275 ;
        RECT 114.570 206.075 115.760 206.360 ;
        RECT 118.690 205.955 120.000 206.275 ;
        RECT 124.370 205.970 124.750 206.350 ;
        RECT 130.030 206.075 131.220 206.360 ;
        RECT 11.820 205.510 12.200 205.890 ;
        RECT 18.275 205.540 18.655 205.920 ;
        RECT 27.280 205.510 27.660 205.890 ;
        RECT 31.025 205.550 31.405 205.930 ;
        RECT 33.735 205.540 34.115 205.920 ;
        RECT 35.145 205.385 38.325 205.705 ;
        RECT 110.045 205.370 110.425 205.750 ;
        RECT 113.790 205.410 114.170 205.790 ;
        RECT 116.500 205.400 116.880 205.780 ;
        RECT 44.650 204.940 45.935 205.320 ;
        RECT 63.965 204.940 65.450 205.320 ;
        RECT 117.910 205.245 121.090 205.565 ;
        RECT 129.250 205.410 129.630 205.790 ;
        RECT 133.370 205.245 136.550 205.565 ;
        RECT 81.130 204.800 82.620 205.180 ;
        RECT 104.820 204.800 105.895 205.180 ;
        RECT 44.110 204.250 45.200 204.630 ;
        RECT 48.595 204.255 61.445 204.590 ;
        RECT 65.610 204.585 65.990 204.630 ;
        RECT 64.875 204.285 66.185 204.585 ;
        RECT 65.610 204.250 65.990 204.285 ;
        RECT 82.780 204.110 83.870 204.490 ;
        RECT 87.265 204.115 100.115 204.450 ;
        RECT 104.280 204.445 104.660 204.490 ;
        RECT 103.545 204.145 104.855 204.445 ;
        RECT 123.650 204.160 127.800 204.430 ;
        RECT 104.280 204.110 104.660 204.145 ;
        RECT 40.965 203.615 74.045 203.740 ;
        RECT 40.965 203.390 106.290 203.615 ;
        RECT 73.340 203.250 106.290 203.390 ;
        RECT 108.085 203.240 112.345 203.595 ;
        RECT 40.935 196.130 78.485 196.140 ;
        RECT 40.935 195.855 106.615 196.130 ;
        RECT 77.840 195.845 106.615 195.855 ;
        RECT 108.285 195.825 114.990 196.125 ;
        RECT 44.640 194.945 45.840 195.325 ;
        RECT 64.165 195.045 65.400 195.425 ;
        RECT 81.145 194.935 82.600 195.315 ;
        RECT 104.840 195.035 106.120 195.415 ;
        RECT 65.580 194.690 65.960 194.725 ;
        RECT 44.080 194.585 44.460 194.625 ;
        RECT 44.010 194.280 46.845 194.585 ;
        RECT 62.825 194.380 65.960 194.690 ;
        RECT 104.280 194.680 104.660 194.715 ;
        RECT 82.780 194.575 83.160 194.615 ;
        RECT 65.580 194.345 65.960 194.380 ;
        RECT 44.080 194.245 44.460 194.280 ;
        RECT 82.710 194.270 85.545 194.575 ;
        RECT 101.525 194.370 104.660 194.680 ;
        RECT 123.790 194.655 130.530 194.955 ;
        RECT 104.280 194.335 104.660 194.370 ;
        RECT 82.780 194.235 83.160 194.270 ;
        RECT 14.410 192.670 14.790 193.050 ;
        RECT 21.310 192.660 21.690 193.040 ;
        RECT 26.125 192.870 29.530 193.310 ;
        RECT 29.870 192.670 30.250 193.050 ;
        RECT 32.585 192.710 32.965 193.090 ;
        RECT 36.770 192.660 37.150 193.040 ;
        RECT 44.640 192.645 47.900 193.025 ;
        RECT 48.640 192.645 51.900 193.025 ;
        RECT 58.140 192.645 61.400 193.025 ;
        RECT 62.140 192.645 65.400 193.025 ;
        RECT 11.735 192.245 13.475 192.535 ;
        RECT 18.235 192.165 20.845 192.590 ;
        RECT 27.195 192.245 28.935 192.535 ;
        RECT 30.985 192.195 32.185 192.485 ;
        RECT 33.695 192.165 36.290 192.540 ;
        RECT 37.905 192.260 38.285 192.640 ;
        RECT 81.305 192.635 82.600 193.015 ;
        RECT 87.340 192.635 90.600 193.015 ;
        RECT 91.340 192.635 92.525 193.015 ;
        RECT 94.790 192.635 96.100 193.015 ;
        RECT 96.840 192.635 100.100 193.015 ;
        RECT 104.840 192.635 105.855 193.015 ;
        RECT 108.920 192.880 112.335 193.300 ;
        RECT 112.665 192.660 113.045 193.040 ;
        RECT 115.380 192.700 115.760 193.080 ;
        RECT 119.565 192.650 119.945 193.030 ;
        RECT 124.380 192.860 127.835 193.300 ;
        RECT 130.840 192.700 131.220 193.080 ;
        RECT 44.080 191.945 44.460 192.325 ;
        RECT 48.080 191.945 48.460 192.325 ;
        RECT 52.080 192.280 52.460 192.325 ;
        RECT 57.580 192.280 57.960 192.325 ;
        RECT 52.030 191.965 57.965 192.280 ;
        RECT 52.080 191.945 52.460 191.965 ;
        RECT 57.580 191.945 57.960 191.965 ;
        RECT 61.580 191.945 61.960 192.325 ;
        RECT 65.580 191.945 65.960 192.325 ;
        RECT 82.780 191.935 83.160 192.315 ;
        RECT 86.780 191.935 87.160 192.315 ;
        RECT 90.780 192.270 91.160 192.315 ;
        RECT 96.280 192.270 96.660 192.315 ;
        RECT 90.730 191.955 96.665 192.270 ;
        RECT 90.780 191.935 91.160 191.955 ;
        RECT 96.280 191.935 96.660 191.955 ;
        RECT 100.280 191.935 100.660 192.315 ;
        RECT 104.280 191.935 104.660 192.315 ;
        RECT 109.990 192.235 111.730 192.525 ;
        RECT 113.780 192.185 114.980 192.475 ;
        RECT 116.490 192.145 119.120 192.600 ;
        RECT 120.700 192.250 121.080 192.630 ;
        RECT 129.240 192.185 130.440 192.475 ;
        RECT 136.160 192.250 136.540 192.630 ;
        RECT 74.870 191.310 95.645 191.685 ;
        RECT 123.195 191.475 139.115 191.775 ;
        RECT 45.305 190.730 72.615 191.070 ;
        RECT 123.730 190.730 140.675 191.030 ;
        RECT 24.920 190.025 32.180 190.325 ;
        RECT 20.420 189.725 23.525 190.000 ;
        RECT 25.475 189.490 29.560 189.760 ;
        RECT 35.880 189.725 39.630 190.000 ;
        RECT 73.900 189.955 105.865 190.345 ;
        RECT 118.675 189.715 121.805 189.990 ;
        RECT 40.935 189.600 59.605 189.610 ;
        RECT 40.935 189.590 98.305 189.600 ;
        RECT 40.935 189.290 107.310 189.590 ;
        RECT 70.745 189.280 107.310 189.290 ;
        RECT 124.925 188.820 129.055 189.120 ;
        RECT 131.430 188.770 135.930 189.080 ;
        RECT 40.405 188.610 76.315 188.620 ;
        RECT 29.135 188.230 35.525 188.520 ;
        RECT 40.405 188.350 107.710 188.610 ;
        RECT 75.965 188.340 107.710 188.350 ;
        RECT 111.930 188.220 118.320 188.510 ;
        RECT 127.390 188.220 133.780 188.510 ;
        RECT 13.090 187.650 23.745 187.985 ;
        RECT 28.550 187.650 39.055 187.985 ;
        RECT 64.025 187.785 74.575 188.120 ;
        RECT 111.345 187.640 121.825 187.975 ;
        RECT 44.620 187.145 47.920 187.525 ;
        RECT 48.620 187.145 51.920 187.525 ;
        RECT 58.120 187.145 61.420 187.525 ;
        RECT 62.120 187.145 65.420 187.525 ;
        RECT 81.315 187.135 82.620 187.515 ;
        RECT 87.320 187.135 90.620 187.515 ;
        RECT 91.320 187.135 92.680 187.515 ;
        RECT 94.655 187.135 96.120 187.515 ;
        RECT 96.820 187.135 100.120 187.515 ;
        RECT 104.820 187.135 106.000 187.515 ;
        RECT 126.155 187.055 129.075 187.355 ;
        RECT 132.620 187.040 135.990 187.340 ;
        RECT 44.080 186.800 44.460 186.835 ;
        RECT 13.060 186.330 14.840 186.620 ;
        RECT 20.435 186.300 21.745 186.620 ;
        RECT 26.115 186.315 26.495 186.695 ;
        RECT 28.520 186.330 30.300 186.620 ;
        RECT 31.775 186.420 32.965 186.705 ;
        RECT 35.895 186.300 37.205 186.620 ;
        RECT 43.815 186.490 46.825 186.800 ;
        RECT 44.080 186.455 44.460 186.490 ;
        RECT 48.080 186.455 49.170 186.835 ;
        RECT 52.080 186.830 52.460 186.835 ;
        RECT 49.600 186.465 52.465 186.830 ;
        RECT 57.580 186.810 57.960 186.835 ;
        RECT 57.565 186.490 59.710 186.810 ;
        RECT 52.080 186.455 52.460 186.465 ;
        RECT 57.580 186.455 57.960 186.490 ;
        RECT 60.625 186.455 61.960 186.835 ;
        RECT 65.580 186.815 65.960 186.835 ;
        RECT 63.115 186.495 66.025 186.815 ;
        RECT 82.780 186.790 83.160 186.825 ;
        RECT 65.580 186.455 65.960 186.495 ;
        RECT 82.515 186.480 85.525 186.790 ;
        RECT 82.780 186.445 83.160 186.480 ;
        RECT 86.780 186.445 87.870 186.825 ;
        RECT 90.780 186.820 91.160 186.825 ;
        RECT 88.300 186.455 91.165 186.820 ;
        RECT 96.280 186.800 96.660 186.825 ;
        RECT 96.265 186.480 98.410 186.800 ;
        RECT 90.780 186.445 91.160 186.455 ;
        RECT 96.280 186.445 96.660 186.480 ;
        RECT 99.325 186.445 100.660 186.825 ;
        RECT 104.280 186.805 104.660 186.825 ;
        RECT 101.815 186.485 104.725 186.805 ;
        RECT 104.280 186.445 104.660 186.485 ;
        RECT 108.910 186.305 109.290 186.685 ;
        RECT 111.315 186.320 113.095 186.610 ;
        RECT 114.570 186.410 115.760 186.695 ;
        RECT 118.690 186.290 120.000 186.610 ;
        RECT 124.370 186.305 124.750 186.685 ;
        RECT 130.030 186.410 131.220 186.695 ;
        RECT 11.790 185.715 12.170 186.095 ;
        RECT 18.245 185.745 18.625 186.125 ;
        RECT 27.250 185.715 27.630 186.095 ;
        RECT 30.995 185.755 31.375 186.135 ;
        RECT 33.705 185.745 34.085 186.125 ;
        RECT 35.115 185.590 38.295 185.910 ;
        RECT 110.045 185.705 110.425 186.085 ;
        RECT 113.790 185.745 114.170 186.125 ;
        RECT 116.500 185.735 116.880 186.115 ;
        RECT 117.910 185.580 121.090 185.900 ;
        RECT 129.250 185.745 129.630 186.125 ;
        RECT 133.370 185.580 136.550 185.900 ;
        RECT 44.620 185.145 45.905 185.525 ;
        RECT 63.935 185.145 65.420 185.525 ;
        RECT 81.130 185.135 82.620 185.515 ;
        RECT 104.820 185.135 105.895 185.515 ;
        RECT 44.080 184.455 45.170 184.835 ;
        RECT 48.565 184.460 61.415 184.795 ;
        RECT 65.580 184.790 65.960 184.835 ;
        RECT 64.845 184.490 66.155 184.790 ;
        RECT 65.580 184.455 65.960 184.490 ;
        RECT 82.780 184.445 83.870 184.825 ;
        RECT 87.265 184.450 100.115 184.785 ;
        RECT 104.280 184.780 104.660 184.825 ;
        RECT 103.545 184.480 104.855 184.780 ;
        RECT 123.650 184.495 127.800 184.765 ;
        RECT 104.280 184.445 104.660 184.480 ;
        RECT 73.340 183.945 106.290 183.950 ;
        RECT 40.935 183.595 106.290 183.945 ;
        RECT 73.340 183.585 106.290 183.595 ;
        RECT 108.085 183.575 112.345 183.930 ;
        RECT 41.085 176.290 78.635 176.345 ;
        RECT 41.085 176.060 106.655 176.290 ;
        RECT 77.880 176.005 106.655 176.060 ;
        RECT 108.325 175.985 115.030 176.285 ;
        RECT 44.790 175.150 45.990 175.530 ;
        RECT 64.315 175.250 65.550 175.630 ;
        RECT 81.185 175.095 82.640 175.475 ;
        RECT 104.880 175.195 106.160 175.575 ;
        RECT 65.730 174.895 66.110 174.930 ;
        RECT 44.230 174.790 44.610 174.830 ;
        RECT 44.160 174.485 46.995 174.790 ;
        RECT 62.975 174.585 66.110 174.895 ;
        RECT 104.320 174.840 104.700 174.875 ;
        RECT 82.820 174.735 83.200 174.775 ;
        RECT 65.730 174.550 66.110 174.585 ;
        RECT 44.230 174.450 44.610 174.485 ;
        RECT 82.750 174.430 85.585 174.735 ;
        RECT 101.565 174.530 104.700 174.840 ;
        RECT 123.830 174.815 130.570 175.115 ;
        RECT 104.320 174.495 104.700 174.530 ;
        RECT 82.820 174.395 83.200 174.430 ;
        RECT 14.560 172.875 14.940 173.255 ;
        RECT 21.460 172.865 21.840 173.245 ;
        RECT 26.275 173.075 29.680 173.515 ;
        RECT 30.020 172.875 30.400 173.255 ;
        RECT 32.735 172.915 33.115 173.295 ;
        RECT 36.920 172.865 37.300 173.245 ;
        RECT 44.790 172.850 48.050 173.230 ;
        RECT 48.790 172.850 52.050 173.230 ;
        RECT 58.290 172.850 61.550 173.230 ;
        RECT 62.290 172.850 65.550 173.230 ;
        RECT 11.885 172.450 13.625 172.740 ;
        RECT 18.385 172.370 20.995 172.795 ;
        RECT 27.345 172.450 29.085 172.740 ;
        RECT 31.135 172.400 32.335 172.690 ;
        RECT 33.845 172.370 36.440 172.745 ;
        RECT 38.055 172.465 38.435 172.845 ;
        RECT 81.345 172.795 82.640 173.175 ;
        RECT 87.380 172.795 90.640 173.175 ;
        RECT 91.380 172.795 92.565 173.175 ;
        RECT 94.830 172.795 96.140 173.175 ;
        RECT 96.880 172.795 100.140 173.175 ;
        RECT 104.880 172.795 105.895 173.175 ;
        RECT 108.960 173.040 112.375 173.460 ;
        RECT 112.705 172.820 113.085 173.200 ;
        RECT 115.420 172.860 115.800 173.240 ;
        RECT 119.605 172.810 119.985 173.190 ;
        RECT 124.420 173.020 127.875 173.460 ;
        RECT 130.880 172.860 131.260 173.240 ;
        RECT 44.230 172.150 44.610 172.530 ;
        RECT 48.230 172.150 48.610 172.530 ;
        RECT 52.230 172.485 52.610 172.530 ;
        RECT 57.730 172.485 58.110 172.530 ;
        RECT 52.180 172.170 58.115 172.485 ;
        RECT 52.230 172.150 52.610 172.170 ;
        RECT 57.730 172.150 58.110 172.170 ;
        RECT 61.730 172.150 62.110 172.530 ;
        RECT 65.730 172.150 66.110 172.530 ;
        RECT 82.820 172.095 83.200 172.475 ;
        RECT 86.820 172.095 87.200 172.475 ;
        RECT 90.820 172.430 91.200 172.475 ;
        RECT 96.320 172.430 96.700 172.475 ;
        RECT 90.770 172.115 96.705 172.430 ;
        RECT 90.820 172.095 91.200 172.115 ;
        RECT 96.320 172.095 96.700 172.115 ;
        RECT 100.320 172.095 100.700 172.475 ;
        RECT 104.320 172.095 104.700 172.475 ;
        RECT 110.030 172.395 111.770 172.685 ;
        RECT 113.820 172.345 115.020 172.635 ;
        RECT 116.530 172.305 119.160 172.760 ;
        RECT 120.740 172.410 121.120 172.790 ;
        RECT 129.280 172.345 130.480 172.635 ;
        RECT 136.200 172.410 136.580 172.790 ;
        RECT 74.910 171.470 95.685 171.845 ;
        RECT 123.235 171.635 139.155 171.935 ;
        RECT 45.455 170.935 72.765 171.275 ;
        RECT 123.770 170.890 140.715 171.190 ;
        RECT 25.070 170.230 32.330 170.530 ;
        RECT 20.570 169.930 23.675 170.205 ;
        RECT 25.625 169.695 29.710 169.965 ;
        RECT 36.030 169.930 39.780 170.205 ;
        RECT 73.940 170.115 105.905 170.505 ;
        RECT 118.715 169.875 121.845 170.150 ;
        RECT 41.085 169.805 59.755 169.815 ;
        RECT 41.085 169.760 71.105 169.805 ;
        RECT 41.085 169.750 98.345 169.760 ;
        RECT 41.085 169.495 107.350 169.750 ;
        RECT 70.785 169.440 107.350 169.495 ;
        RECT 124.965 168.980 129.095 169.280 ;
        RECT 131.470 168.930 135.970 169.240 ;
        RECT 40.555 168.770 76.465 168.825 ;
        RECT 29.285 168.435 35.675 168.725 ;
        RECT 40.555 168.555 107.750 168.770 ;
        RECT 76.005 168.500 107.750 168.555 ;
        RECT 111.970 168.380 118.360 168.670 ;
        RECT 127.430 168.380 133.820 168.670 ;
        RECT 13.240 167.855 23.895 168.190 ;
        RECT 28.700 167.855 39.205 168.190 ;
        RECT 64.175 167.990 74.725 168.325 ;
        RECT 111.385 167.800 121.865 168.135 ;
        RECT 44.770 167.350 48.070 167.730 ;
        RECT 48.770 167.350 52.070 167.730 ;
        RECT 58.270 167.350 61.570 167.730 ;
        RECT 62.270 167.350 65.570 167.730 ;
        RECT 81.355 167.295 82.660 167.675 ;
        RECT 87.360 167.295 90.660 167.675 ;
        RECT 91.360 167.295 92.720 167.675 ;
        RECT 94.695 167.295 96.160 167.675 ;
        RECT 96.860 167.295 100.160 167.675 ;
        RECT 104.860 167.295 106.040 167.675 ;
        RECT 126.195 167.215 129.115 167.515 ;
        RECT 132.660 167.200 136.030 167.500 ;
        RECT 44.230 167.005 44.610 167.040 ;
        RECT 13.210 166.535 14.990 166.825 ;
        RECT 20.585 166.505 21.895 166.825 ;
        RECT 26.265 166.520 26.645 166.900 ;
        RECT 28.670 166.535 30.450 166.825 ;
        RECT 31.925 166.625 33.115 166.910 ;
        RECT 36.045 166.505 37.355 166.825 ;
        RECT 43.965 166.695 46.975 167.005 ;
        RECT 44.230 166.660 44.610 166.695 ;
        RECT 48.230 166.660 49.320 167.040 ;
        RECT 52.230 167.035 52.610 167.040 ;
        RECT 49.750 166.670 52.615 167.035 ;
        RECT 57.730 167.015 58.110 167.040 ;
        RECT 57.715 166.695 59.860 167.015 ;
        RECT 52.230 166.660 52.610 166.670 ;
        RECT 57.730 166.660 58.110 166.695 ;
        RECT 60.775 166.660 62.110 167.040 ;
        RECT 65.730 167.020 66.110 167.040 ;
        RECT 63.265 166.700 66.175 167.020 ;
        RECT 82.820 166.950 83.200 166.985 ;
        RECT 65.730 166.660 66.110 166.700 ;
        RECT 82.555 166.640 85.565 166.950 ;
        RECT 82.820 166.605 83.200 166.640 ;
        RECT 86.820 166.605 87.910 166.985 ;
        RECT 90.820 166.980 91.200 166.985 ;
        RECT 88.340 166.615 91.205 166.980 ;
        RECT 96.320 166.960 96.700 166.985 ;
        RECT 96.305 166.640 98.450 166.960 ;
        RECT 90.820 166.605 91.200 166.615 ;
        RECT 96.320 166.605 96.700 166.640 ;
        RECT 99.365 166.605 100.700 166.985 ;
        RECT 104.320 166.965 104.700 166.985 ;
        RECT 101.855 166.645 104.765 166.965 ;
        RECT 104.320 166.605 104.700 166.645 ;
        RECT 108.950 166.465 109.330 166.845 ;
        RECT 111.355 166.480 113.135 166.770 ;
        RECT 114.610 166.570 115.800 166.855 ;
        RECT 118.730 166.450 120.040 166.770 ;
        RECT 124.410 166.465 124.790 166.845 ;
        RECT 130.070 166.570 131.260 166.855 ;
        RECT 11.940 165.920 12.320 166.300 ;
        RECT 18.395 165.950 18.775 166.330 ;
        RECT 27.400 165.920 27.780 166.300 ;
        RECT 31.145 165.960 31.525 166.340 ;
        RECT 33.855 165.950 34.235 166.330 ;
        RECT 35.265 165.795 38.445 166.115 ;
        RECT 110.085 165.865 110.465 166.245 ;
        RECT 113.830 165.905 114.210 166.285 ;
        RECT 116.540 165.895 116.920 166.275 ;
        RECT 117.950 165.740 121.130 166.060 ;
        RECT 129.290 165.905 129.670 166.285 ;
        RECT 133.410 165.740 136.590 166.060 ;
        RECT 44.770 165.350 46.055 165.730 ;
        RECT 64.085 165.350 65.570 165.730 ;
        RECT 81.170 165.295 82.660 165.675 ;
        RECT 104.860 165.295 105.935 165.675 ;
        RECT 44.230 164.660 45.320 165.040 ;
        RECT 48.715 164.665 61.565 165.000 ;
        RECT 65.730 164.995 66.110 165.040 ;
        RECT 64.995 164.695 66.305 164.995 ;
        RECT 65.730 164.660 66.110 164.695 ;
        RECT 82.820 164.605 83.910 164.985 ;
        RECT 87.305 164.610 100.155 164.945 ;
        RECT 104.320 164.940 104.700 164.985 ;
        RECT 103.585 164.640 104.895 164.940 ;
        RECT 123.690 164.655 127.840 164.925 ;
        RECT 104.320 164.605 104.700 164.640 ;
        RECT 41.085 164.110 74.165 164.150 ;
        RECT 41.085 163.800 106.330 164.110 ;
        RECT 73.380 163.745 106.330 163.800 ;
        RECT 108.125 163.735 112.385 164.090 ;
        RECT 41.040 156.565 78.590 156.655 ;
        RECT 41.040 156.370 106.455 156.565 ;
        RECT 77.680 156.280 106.455 156.370 ;
        RECT 108.125 156.260 114.830 156.560 ;
        RECT 44.745 155.460 45.945 155.840 ;
        RECT 64.270 155.560 65.505 155.940 ;
        RECT 80.985 155.370 82.440 155.750 ;
        RECT 104.680 155.470 105.960 155.850 ;
        RECT 65.685 155.205 66.065 155.240 ;
        RECT 44.185 155.100 44.565 155.140 ;
        RECT 44.115 154.795 46.950 155.100 ;
        RECT 62.930 154.895 66.065 155.205 ;
        RECT 104.120 155.115 104.500 155.150 ;
        RECT 82.620 155.010 83.000 155.050 ;
        RECT 65.685 154.860 66.065 154.895 ;
        RECT 44.185 154.760 44.565 154.795 ;
        RECT 82.550 154.705 85.385 155.010 ;
        RECT 101.365 154.805 104.500 155.115 ;
        RECT 123.630 155.090 130.370 155.390 ;
        RECT 104.120 154.770 104.500 154.805 ;
        RECT 82.620 154.670 83.000 154.705 ;
        RECT 14.515 153.185 14.895 153.565 ;
        RECT 21.415 153.175 21.795 153.555 ;
        RECT 26.230 153.385 29.635 153.825 ;
        RECT 29.975 153.185 30.355 153.565 ;
        RECT 32.690 153.225 33.070 153.605 ;
        RECT 36.875 153.175 37.255 153.555 ;
        RECT 44.745 153.160 48.005 153.540 ;
        RECT 48.745 153.160 52.005 153.540 ;
        RECT 58.245 153.160 61.505 153.540 ;
        RECT 62.245 153.160 65.505 153.540 ;
        RECT 11.840 152.760 13.580 153.050 ;
        RECT 18.340 152.680 20.950 153.105 ;
        RECT 27.300 152.760 29.040 153.050 ;
        RECT 31.090 152.710 32.290 153.000 ;
        RECT 33.800 152.680 36.395 153.055 ;
        RECT 38.010 152.775 38.390 153.155 ;
        RECT 81.145 153.070 82.440 153.450 ;
        RECT 87.180 153.070 90.440 153.450 ;
        RECT 91.180 153.070 92.365 153.450 ;
        RECT 94.630 153.070 95.940 153.450 ;
        RECT 96.680 153.070 99.940 153.450 ;
        RECT 104.680 153.070 105.695 153.450 ;
        RECT 108.760 153.315 112.175 153.735 ;
        RECT 112.505 153.095 112.885 153.475 ;
        RECT 115.220 153.135 115.600 153.515 ;
        RECT 119.405 153.085 119.785 153.465 ;
        RECT 124.220 153.295 127.675 153.735 ;
        RECT 130.680 153.135 131.060 153.515 ;
        RECT 44.185 152.460 44.565 152.840 ;
        RECT 48.185 152.460 48.565 152.840 ;
        RECT 52.185 152.795 52.565 152.840 ;
        RECT 57.685 152.795 58.065 152.840 ;
        RECT 52.135 152.480 58.070 152.795 ;
        RECT 52.185 152.460 52.565 152.480 ;
        RECT 57.685 152.460 58.065 152.480 ;
        RECT 61.685 152.460 62.065 152.840 ;
        RECT 65.685 152.460 66.065 152.840 ;
        RECT 82.620 152.370 83.000 152.750 ;
        RECT 86.620 152.370 87.000 152.750 ;
        RECT 90.620 152.705 91.000 152.750 ;
        RECT 96.120 152.705 96.500 152.750 ;
        RECT 90.570 152.390 96.505 152.705 ;
        RECT 90.620 152.370 91.000 152.390 ;
        RECT 96.120 152.370 96.500 152.390 ;
        RECT 100.120 152.370 100.500 152.750 ;
        RECT 104.120 152.370 104.500 152.750 ;
        RECT 109.830 152.670 111.570 152.960 ;
        RECT 113.620 152.620 114.820 152.910 ;
        RECT 116.330 152.580 118.960 153.035 ;
        RECT 120.540 152.685 120.920 153.065 ;
        RECT 129.080 152.620 130.280 152.910 ;
        RECT 136.000 152.685 136.380 153.065 ;
        RECT 74.710 151.745 95.485 152.120 ;
        RECT 123.035 151.910 138.955 152.210 ;
        RECT 45.410 151.245 72.720 151.585 ;
        RECT 123.570 151.165 140.515 151.465 ;
        RECT 25.025 150.540 32.285 150.840 ;
        RECT 20.525 150.240 23.630 150.515 ;
        RECT 25.580 150.005 29.665 150.275 ;
        RECT 35.985 150.240 39.735 150.515 ;
        RECT 73.740 150.390 105.705 150.780 ;
        RECT 118.515 150.150 121.645 150.425 ;
        RECT 41.040 150.115 59.710 150.125 ;
        RECT 41.040 150.035 71.060 150.115 ;
        RECT 41.040 150.025 98.145 150.035 ;
        RECT 41.040 149.805 107.150 150.025 ;
        RECT 70.585 149.715 107.150 149.805 ;
        RECT 124.765 149.255 128.895 149.555 ;
        RECT 131.270 149.205 135.770 149.515 ;
        RECT 40.510 149.045 76.420 149.135 ;
        RECT 29.240 148.745 35.630 149.035 ;
        RECT 40.510 148.865 107.550 149.045 ;
        RECT 75.805 148.775 107.550 148.865 ;
        RECT 111.770 148.655 118.160 148.945 ;
        RECT 127.230 148.655 133.620 148.945 ;
        RECT 13.195 148.165 23.850 148.500 ;
        RECT 28.655 148.165 39.160 148.500 ;
        RECT 64.130 148.300 74.680 148.635 ;
        RECT 111.185 148.075 121.665 148.410 ;
        RECT 44.725 147.660 48.025 148.040 ;
        RECT 48.725 147.660 52.025 148.040 ;
        RECT 58.225 147.660 61.525 148.040 ;
        RECT 62.225 147.660 65.525 148.040 ;
        RECT 81.155 147.570 82.460 147.950 ;
        RECT 87.160 147.570 90.460 147.950 ;
        RECT 91.160 147.570 92.520 147.950 ;
        RECT 94.495 147.570 95.960 147.950 ;
        RECT 96.660 147.570 99.960 147.950 ;
        RECT 104.660 147.570 105.840 147.950 ;
        RECT 125.995 147.490 128.915 147.790 ;
        RECT 132.460 147.475 135.830 147.775 ;
        RECT 44.185 147.315 44.565 147.350 ;
        RECT 13.165 146.845 14.945 147.135 ;
        RECT 20.540 146.815 21.850 147.135 ;
        RECT 26.220 146.830 26.600 147.210 ;
        RECT 28.625 146.845 30.405 147.135 ;
        RECT 31.880 146.935 33.070 147.220 ;
        RECT 36.000 146.815 37.310 147.135 ;
        RECT 43.920 147.005 46.930 147.315 ;
        RECT 44.185 146.970 44.565 147.005 ;
        RECT 48.185 146.970 49.275 147.350 ;
        RECT 52.185 147.345 52.565 147.350 ;
        RECT 49.705 146.980 52.570 147.345 ;
        RECT 57.685 147.325 58.065 147.350 ;
        RECT 57.670 147.005 59.815 147.325 ;
        RECT 52.185 146.970 52.565 146.980 ;
        RECT 57.685 146.970 58.065 147.005 ;
        RECT 60.730 146.970 62.065 147.350 ;
        RECT 65.685 147.330 66.065 147.350 ;
        RECT 63.220 147.010 66.130 147.330 ;
        RECT 82.620 147.225 83.000 147.260 ;
        RECT 65.685 146.970 66.065 147.010 ;
        RECT 82.355 146.915 85.365 147.225 ;
        RECT 82.620 146.880 83.000 146.915 ;
        RECT 86.620 146.880 87.710 147.260 ;
        RECT 90.620 147.255 91.000 147.260 ;
        RECT 88.140 146.890 91.005 147.255 ;
        RECT 96.120 147.235 96.500 147.260 ;
        RECT 96.105 146.915 98.250 147.235 ;
        RECT 90.620 146.880 91.000 146.890 ;
        RECT 96.120 146.880 96.500 146.915 ;
        RECT 99.165 146.880 100.500 147.260 ;
        RECT 104.120 147.240 104.500 147.260 ;
        RECT 101.655 146.920 104.565 147.240 ;
        RECT 104.120 146.880 104.500 146.920 ;
        RECT 108.750 146.740 109.130 147.120 ;
        RECT 111.155 146.755 112.935 147.045 ;
        RECT 114.410 146.845 115.600 147.130 ;
        RECT 118.530 146.725 119.840 147.045 ;
        RECT 124.210 146.740 124.590 147.120 ;
        RECT 129.870 146.845 131.060 147.130 ;
        RECT 11.895 146.230 12.275 146.610 ;
        RECT 18.350 146.260 18.730 146.640 ;
        RECT 27.355 146.230 27.735 146.610 ;
        RECT 31.100 146.270 31.480 146.650 ;
        RECT 33.810 146.260 34.190 146.640 ;
        RECT 35.220 146.105 38.400 146.425 ;
        RECT 109.885 146.140 110.265 146.520 ;
        RECT 113.630 146.180 114.010 146.560 ;
        RECT 116.340 146.170 116.720 146.550 ;
        RECT 44.725 145.660 46.010 146.040 ;
        RECT 64.040 145.660 65.525 146.040 ;
        RECT 117.750 146.015 120.930 146.335 ;
        RECT 129.090 146.180 129.470 146.560 ;
        RECT 133.210 146.015 136.390 146.335 ;
        RECT 80.970 145.570 82.460 145.950 ;
        RECT 104.660 145.570 105.735 145.950 ;
        RECT 44.185 144.970 45.275 145.350 ;
        RECT 48.670 144.975 61.520 145.310 ;
        RECT 65.685 145.305 66.065 145.350 ;
        RECT 64.950 145.005 66.260 145.305 ;
        RECT 65.685 144.970 66.065 145.005 ;
        RECT 82.620 144.880 83.710 145.260 ;
        RECT 87.105 144.885 99.955 145.220 ;
        RECT 104.120 145.215 104.500 145.260 ;
        RECT 103.385 144.915 104.695 145.215 ;
        RECT 123.490 144.930 127.640 145.200 ;
        RECT 104.120 144.880 104.500 144.915 ;
        RECT 41.040 144.385 74.120 144.460 ;
        RECT 41.040 144.110 106.130 144.385 ;
        RECT 73.180 144.020 106.130 144.110 ;
        RECT 107.925 144.010 112.185 144.365 ;
        RECT 41.230 136.920 78.780 136.945 ;
        RECT 41.230 136.660 106.610 136.920 ;
        RECT 77.835 136.635 106.610 136.660 ;
        RECT 108.280 136.615 114.985 136.915 ;
        RECT 44.935 135.750 46.135 136.130 ;
        RECT 64.460 135.850 65.695 136.230 ;
        RECT 81.140 135.725 82.595 136.105 ;
        RECT 104.835 135.825 106.115 136.205 ;
        RECT 65.875 135.495 66.255 135.530 ;
        RECT 44.375 135.390 44.755 135.430 ;
        RECT 44.305 135.085 47.140 135.390 ;
        RECT 63.120 135.185 66.255 135.495 ;
        RECT 104.275 135.470 104.655 135.505 ;
        RECT 82.775 135.365 83.155 135.405 ;
        RECT 65.875 135.150 66.255 135.185 ;
        RECT 44.375 135.050 44.755 135.085 ;
        RECT 82.705 135.060 85.540 135.365 ;
        RECT 101.520 135.160 104.655 135.470 ;
        RECT 123.785 135.445 130.525 135.745 ;
        RECT 104.275 135.125 104.655 135.160 ;
        RECT 82.775 135.025 83.155 135.060 ;
        RECT 14.705 133.475 15.085 133.855 ;
        RECT 21.605 133.465 21.985 133.845 ;
        RECT 26.420 133.675 29.825 134.115 ;
        RECT 30.165 133.475 30.545 133.855 ;
        RECT 32.880 133.515 33.260 133.895 ;
        RECT 37.065 133.465 37.445 133.845 ;
        RECT 44.935 133.450 48.195 133.830 ;
        RECT 48.935 133.450 52.195 133.830 ;
        RECT 58.435 133.450 61.695 133.830 ;
        RECT 62.435 133.450 65.695 133.830 ;
        RECT 12.030 133.050 13.770 133.340 ;
        RECT 18.530 132.970 21.140 133.395 ;
        RECT 27.490 133.050 29.230 133.340 ;
        RECT 31.280 133.000 32.480 133.290 ;
        RECT 33.990 132.970 36.585 133.345 ;
        RECT 38.200 133.065 38.580 133.445 ;
        RECT 81.300 133.425 82.595 133.805 ;
        RECT 87.335 133.425 90.595 133.805 ;
        RECT 91.335 133.425 92.520 133.805 ;
        RECT 94.785 133.425 96.095 133.805 ;
        RECT 96.835 133.425 100.095 133.805 ;
        RECT 104.835 133.425 105.850 133.805 ;
        RECT 108.915 133.670 112.330 134.090 ;
        RECT 112.660 133.450 113.040 133.830 ;
        RECT 115.375 133.490 115.755 133.870 ;
        RECT 119.560 133.440 119.940 133.820 ;
        RECT 124.375 133.650 127.830 134.090 ;
        RECT 130.835 133.490 131.215 133.870 ;
        RECT 44.375 132.750 44.755 133.130 ;
        RECT 48.375 132.750 48.755 133.130 ;
        RECT 52.375 133.085 52.755 133.130 ;
        RECT 57.875 133.085 58.255 133.130 ;
        RECT 52.325 132.770 58.260 133.085 ;
        RECT 52.375 132.750 52.755 132.770 ;
        RECT 57.875 132.750 58.255 132.770 ;
        RECT 61.875 132.750 62.255 133.130 ;
        RECT 65.875 132.750 66.255 133.130 ;
        RECT 82.775 132.725 83.155 133.105 ;
        RECT 86.775 132.725 87.155 133.105 ;
        RECT 90.775 133.060 91.155 133.105 ;
        RECT 96.275 133.060 96.655 133.105 ;
        RECT 90.725 132.745 96.660 133.060 ;
        RECT 90.775 132.725 91.155 132.745 ;
        RECT 96.275 132.725 96.655 132.745 ;
        RECT 100.275 132.725 100.655 133.105 ;
        RECT 104.275 132.725 104.655 133.105 ;
        RECT 109.985 133.025 111.725 133.315 ;
        RECT 113.775 132.975 114.975 133.265 ;
        RECT 116.485 132.935 119.115 133.390 ;
        RECT 120.695 133.040 121.075 133.420 ;
        RECT 129.235 132.975 130.435 133.265 ;
        RECT 136.155 133.040 136.535 133.420 ;
        RECT 74.865 132.100 95.640 132.475 ;
        RECT 123.190 132.265 139.110 132.565 ;
        RECT 45.600 131.535 72.910 131.875 ;
        RECT 123.725 131.520 140.670 131.820 ;
        RECT 25.215 130.830 32.475 131.130 ;
        RECT 20.715 130.530 23.820 130.805 ;
        RECT 25.770 130.295 29.855 130.565 ;
        RECT 36.175 130.530 39.925 130.805 ;
        RECT 73.895 130.745 105.860 131.135 ;
        RECT 118.670 130.505 121.800 130.780 ;
        RECT 41.230 130.405 59.900 130.415 ;
        RECT 41.230 130.390 71.250 130.405 ;
        RECT 41.230 130.380 98.300 130.390 ;
        RECT 41.230 130.095 107.305 130.380 ;
        RECT 70.740 130.070 107.305 130.095 ;
        RECT 124.920 129.610 129.050 129.910 ;
        RECT 131.425 129.560 135.925 129.870 ;
        RECT 40.700 129.400 76.610 129.425 ;
        RECT 29.430 129.035 35.820 129.325 ;
        RECT 40.700 129.155 107.705 129.400 ;
        RECT 75.960 129.130 107.705 129.155 ;
        RECT 111.925 129.010 118.315 129.300 ;
        RECT 127.385 129.010 133.775 129.300 ;
        RECT 13.385 128.455 24.040 128.790 ;
        RECT 28.845 128.455 39.350 128.790 ;
        RECT 64.320 128.590 74.870 128.925 ;
        RECT 111.340 128.430 121.820 128.765 ;
        RECT 44.915 127.950 48.215 128.330 ;
        RECT 48.915 127.950 52.215 128.330 ;
        RECT 58.415 127.950 61.715 128.330 ;
        RECT 62.415 127.950 65.715 128.330 ;
        RECT 81.310 127.925 82.615 128.305 ;
        RECT 87.315 127.925 90.615 128.305 ;
        RECT 91.315 127.925 92.675 128.305 ;
        RECT 94.650 127.925 96.115 128.305 ;
        RECT 96.815 127.925 100.115 128.305 ;
        RECT 104.815 127.925 105.995 128.305 ;
        RECT 126.150 127.845 129.070 128.145 ;
        RECT 132.615 127.830 135.985 128.130 ;
        RECT 44.375 127.605 44.755 127.640 ;
        RECT 13.355 127.135 15.135 127.425 ;
        RECT 20.730 127.105 22.040 127.425 ;
        RECT 26.410 127.120 26.790 127.500 ;
        RECT 28.815 127.135 30.595 127.425 ;
        RECT 32.070 127.225 33.260 127.510 ;
        RECT 36.190 127.105 37.500 127.425 ;
        RECT 44.110 127.295 47.120 127.605 ;
        RECT 44.375 127.260 44.755 127.295 ;
        RECT 48.375 127.260 49.465 127.640 ;
        RECT 52.375 127.635 52.755 127.640 ;
        RECT 49.895 127.270 52.760 127.635 ;
        RECT 57.875 127.615 58.255 127.640 ;
        RECT 57.860 127.295 60.005 127.615 ;
        RECT 52.375 127.260 52.755 127.270 ;
        RECT 57.875 127.260 58.255 127.295 ;
        RECT 60.920 127.260 62.255 127.640 ;
        RECT 65.875 127.620 66.255 127.640 ;
        RECT 63.410 127.300 66.320 127.620 ;
        RECT 82.775 127.580 83.155 127.615 ;
        RECT 65.875 127.260 66.255 127.300 ;
        RECT 82.510 127.270 85.520 127.580 ;
        RECT 82.775 127.235 83.155 127.270 ;
        RECT 86.775 127.235 87.865 127.615 ;
        RECT 90.775 127.610 91.155 127.615 ;
        RECT 88.295 127.245 91.160 127.610 ;
        RECT 96.275 127.590 96.655 127.615 ;
        RECT 96.260 127.270 98.405 127.590 ;
        RECT 90.775 127.235 91.155 127.245 ;
        RECT 96.275 127.235 96.655 127.270 ;
        RECT 99.320 127.235 100.655 127.615 ;
        RECT 104.275 127.595 104.655 127.615 ;
        RECT 101.810 127.275 104.720 127.595 ;
        RECT 104.275 127.235 104.655 127.275 ;
        RECT 108.905 127.095 109.285 127.475 ;
        RECT 111.310 127.110 113.090 127.400 ;
        RECT 114.565 127.200 115.755 127.485 ;
        RECT 118.685 127.080 119.995 127.400 ;
        RECT 124.365 127.095 124.745 127.475 ;
        RECT 130.025 127.200 131.215 127.485 ;
        RECT 12.085 126.520 12.465 126.900 ;
        RECT 18.540 126.550 18.920 126.930 ;
        RECT 27.545 126.520 27.925 126.900 ;
        RECT 31.290 126.560 31.670 126.940 ;
        RECT 34.000 126.550 34.380 126.930 ;
        RECT 35.410 126.395 38.590 126.715 ;
        RECT 110.040 126.495 110.420 126.875 ;
        RECT 113.785 126.535 114.165 126.915 ;
        RECT 116.495 126.525 116.875 126.905 ;
        RECT 117.905 126.370 121.085 126.690 ;
        RECT 129.245 126.535 129.625 126.915 ;
        RECT 133.365 126.370 136.545 126.690 ;
        RECT 44.915 125.950 46.200 126.330 ;
        RECT 64.230 125.950 65.715 126.330 ;
        RECT 81.125 125.925 82.615 126.305 ;
        RECT 104.815 125.925 105.890 126.305 ;
        RECT 44.375 125.260 45.465 125.640 ;
        RECT 48.860 125.265 61.710 125.600 ;
        RECT 65.875 125.595 66.255 125.640 ;
        RECT 65.140 125.295 66.450 125.595 ;
        RECT 65.875 125.260 66.255 125.295 ;
        RECT 82.775 125.235 83.865 125.615 ;
        RECT 87.260 125.240 100.110 125.575 ;
        RECT 104.275 125.570 104.655 125.615 ;
        RECT 103.540 125.270 104.850 125.570 ;
        RECT 123.645 125.285 127.795 125.555 ;
        RECT 104.275 125.235 104.655 125.270 ;
        RECT 41.230 124.740 74.310 124.750 ;
        RECT 41.230 124.400 106.285 124.740 ;
        RECT 73.335 124.375 106.285 124.400 ;
        RECT 108.080 124.365 112.340 124.720 ;
        RECT 77.835 117.105 106.610 117.125 ;
        RECT 41.035 116.840 106.610 117.105 ;
        RECT 41.035 116.820 78.585 116.840 ;
        RECT 108.280 116.820 114.985 117.120 ;
        RECT 44.740 115.910 45.940 116.290 ;
        RECT 64.265 116.010 65.500 116.390 ;
        RECT 81.140 115.930 82.595 116.310 ;
        RECT 104.835 116.030 106.115 116.410 ;
        RECT 65.680 115.655 66.060 115.690 ;
        RECT 104.275 115.675 104.655 115.710 ;
        RECT 44.180 115.550 44.560 115.590 ;
        RECT 44.110 115.245 46.945 115.550 ;
        RECT 62.925 115.345 66.060 115.655 ;
        RECT 82.775 115.570 83.155 115.610 ;
        RECT 65.680 115.310 66.060 115.345 ;
        RECT 82.705 115.265 85.540 115.570 ;
        RECT 101.520 115.365 104.655 115.675 ;
        RECT 123.785 115.650 130.525 115.950 ;
        RECT 104.275 115.330 104.655 115.365 ;
        RECT 44.180 115.210 44.560 115.245 ;
        RECT 82.775 115.230 83.155 115.265 ;
        RECT 14.510 113.635 14.890 114.015 ;
        RECT 21.410 113.625 21.790 114.005 ;
        RECT 26.225 113.835 29.630 114.275 ;
        RECT 29.970 113.635 30.350 114.015 ;
        RECT 32.685 113.675 33.065 114.055 ;
        RECT 36.870 113.625 37.250 114.005 ;
        RECT 44.740 113.610 48.000 113.990 ;
        RECT 48.740 113.610 52.000 113.990 ;
        RECT 58.240 113.610 61.500 113.990 ;
        RECT 62.240 113.610 65.500 113.990 ;
        RECT 81.300 113.630 82.595 114.010 ;
        RECT 87.335 113.630 90.595 114.010 ;
        RECT 91.335 113.630 92.520 114.010 ;
        RECT 94.785 113.630 96.095 114.010 ;
        RECT 96.835 113.630 100.095 114.010 ;
        RECT 104.835 113.630 105.850 114.010 ;
        RECT 108.915 113.875 112.330 114.295 ;
        RECT 112.660 113.655 113.040 114.035 ;
        RECT 115.375 113.695 115.755 114.075 ;
        RECT 119.560 113.645 119.940 114.025 ;
        RECT 124.375 113.855 127.830 114.295 ;
        RECT 130.835 113.695 131.215 114.075 ;
        RECT 11.835 113.210 13.575 113.500 ;
        RECT 18.335 113.130 20.945 113.555 ;
        RECT 27.295 113.210 29.035 113.500 ;
        RECT 31.085 113.160 32.285 113.450 ;
        RECT 33.795 113.130 36.390 113.505 ;
        RECT 38.005 113.225 38.385 113.605 ;
        RECT 44.180 112.910 44.560 113.290 ;
        RECT 48.180 112.910 48.560 113.290 ;
        RECT 52.180 113.245 52.560 113.290 ;
        RECT 57.680 113.245 58.060 113.290 ;
        RECT 52.130 112.930 58.065 113.245 ;
        RECT 52.180 112.910 52.560 112.930 ;
        RECT 57.680 112.910 58.060 112.930 ;
        RECT 61.680 112.910 62.060 113.290 ;
        RECT 65.680 112.910 66.060 113.290 ;
        RECT 82.775 112.930 83.155 113.310 ;
        RECT 86.775 112.930 87.155 113.310 ;
        RECT 90.775 113.265 91.155 113.310 ;
        RECT 96.275 113.265 96.655 113.310 ;
        RECT 90.725 112.950 96.660 113.265 ;
        RECT 90.775 112.930 91.155 112.950 ;
        RECT 96.275 112.930 96.655 112.950 ;
        RECT 100.275 112.930 100.655 113.310 ;
        RECT 104.275 112.930 104.655 113.310 ;
        RECT 109.985 113.230 111.725 113.520 ;
        RECT 113.775 113.180 114.975 113.470 ;
        RECT 116.485 113.140 119.115 113.595 ;
        RECT 120.695 113.245 121.075 113.625 ;
        RECT 129.235 113.180 130.435 113.470 ;
        RECT 136.155 113.245 136.535 113.625 ;
        RECT 74.865 112.305 95.640 112.680 ;
        RECT 123.190 112.470 139.110 112.770 ;
        RECT 45.405 111.695 72.715 112.035 ;
        RECT 123.725 111.725 140.670 112.025 ;
        RECT 25.020 110.990 32.280 111.290 ;
        RECT 20.520 110.690 23.625 110.965 ;
        RECT 25.575 110.455 29.660 110.725 ;
        RECT 35.980 110.690 39.730 110.965 ;
        RECT 73.895 110.950 105.860 111.340 ;
        RECT 118.670 110.710 121.800 110.985 ;
        RECT 70.740 110.585 98.300 110.595 ;
        RECT 41.035 110.565 59.705 110.575 ;
        RECT 70.740 110.565 107.305 110.585 ;
        RECT 41.035 110.275 107.305 110.565 ;
        RECT 41.035 110.255 71.055 110.275 ;
        RECT 124.920 109.815 129.050 110.115 ;
        RECT 131.425 109.765 135.925 110.075 ;
        RECT 75.960 109.585 107.705 109.605 ;
        RECT 29.235 109.195 35.625 109.485 ;
        RECT 40.505 109.335 107.705 109.585 ;
        RECT 40.505 109.315 76.415 109.335 ;
        RECT 111.925 109.215 118.315 109.505 ;
        RECT 127.385 109.215 133.775 109.505 ;
        RECT 13.190 108.615 23.845 108.950 ;
        RECT 28.650 108.615 39.155 108.950 ;
        RECT 64.125 108.750 74.675 109.085 ;
        RECT 111.340 108.635 121.820 108.970 ;
        RECT 44.720 108.110 48.020 108.490 ;
        RECT 48.720 108.110 52.020 108.490 ;
        RECT 58.220 108.110 61.520 108.490 ;
        RECT 62.220 108.110 65.520 108.490 ;
        RECT 81.310 108.130 82.615 108.510 ;
        RECT 87.315 108.130 90.615 108.510 ;
        RECT 91.315 108.130 92.675 108.510 ;
        RECT 94.650 108.130 96.115 108.510 ;
        RECT 96.815 108.130 100.115 108.510 ;
        RECT 104.815 108.130 105.995 108.510 ;
        RECT 126.150 108.050 129.070 108.350 ;
        RECT 132.615 108.035 135.985 108.335 ;
        RECT 44.180 107.765 44.560 107.800 ;
        RECT 13.160 107.295 14.940 107.585 ;
        RECT 20.535 107.265 21.845 107.585 ;
        RECT 26.215 107.280 26.595 107.660 ;
        RECT 28.620 107.295 30.400 107.585 ;
        RECT 31.875 107.385 33.065 107.670 ;
        RECT 35.995 107.265 37.305 107.585 ;
        RECT 43.915 107.455 46.925 107.765 ;
        RECT 44.180 107.420 44.560 107.455 ;
        RECT 48.180 107.420 49.270 107.800 ;
        RECT 52.180 107.795 52.560 107.800 ;
        RECT 49.700 107.430 52.565 107.795 ;
        RECT 57.680 107.775 58.060 107.800 ;
        RECT 57.665 107.455 59.810 107.775 ;
        RECT 52.180 107.420 52.560 107.430 ;
        RECT 57.680 107.420 58.060 107.455 ;
        RECT 60.725 107.420 62.060 107.800 ;
        RECT 65.680 107.780 66.060 107.800 ;
        RECT 82.775 107.785 83.155 107.820 ;
        RECT 63.215 107.460 66.125 107.780 ;
        RECT 82.510 107.475 85.520 107.785 ;
        RECT 65.680 107.420 66.060 107.460 ;
        RECT 82.775 107.440 83.155 107.475 ;
        RECT 86.775 107.440 87.865 107.820 ;
        RECT 90.775 107.815 91.155 107.820 ;
        RECT 88.295 107.450 91.160 107.815 ;
        RECT 96.275 107.795 96.655 107.820 ;
        RECT 96.260 107.475 98.405 107.795 ;
        RECT 90.775 107.440 91.155 107.450 ;
        RECT 96.275 107.440 96.655 107.475 ;
        RECT 99.320 107.440 100.655 107.820 ;
        RECT 104.275 107.800 104.655 107.820 ;
        RECT 101.810 107.480 104.720 107.800 ;
        RECT 104.275 107.440 104.655 107.480 ;
        RECT 108.905 107.300 109.285 107.680 ;
        RECT 111.310 107.315 113.090 107.605 ;
        RECT 114.565 107.405 115.755 107.690 ;
        RECT 118.685 107.285 119.995 107.605 ;
        RECT 124.365 107.300 124.745 107.680 ;
        RECT 130.025 107.405 131.215 107.690 ;
        RECT 11.890 106.680 12.270 107.060 ;
        RECT 18.345 106.710 18.725 107.090 ;
        RECT 27.350 106.680 27.730 107.060 ;
        RECT 31.095 106.720 31.475 107.100 ;
        RECT 33.805 106.710 34.185 107.090 ;
        RECT 35.215 106.555 38.395 106.875 ;
        RECT 110.040 106.700 110.420 107.080 ;
        RECT 113.785 106.740 114.165 107.120 ;
        RECT 116.495 106.730 116.875 107.110 ;
        RECT 117.905 106.575 121.085 106.895 ;
        RECT 129.245 106.740 129.625 107.120 ;
        RECT 133.365 106.575 136.545 106.895 ;
        RECT 44.720 106.110 46.005 106.490 ;
        RECT 64.035 106.110 65.520 106.490 ;
        RECT 81.125 106.130 82.615 106.510 ;
        RECT 104.815 106.130 105.890 106.510 ;
        RECT 44.180 105.420 45.270 105.800 ;
        RECT 48.665 105.425 61.515 105.760 ;
        RECT 65.680 105.755 66.060 105.800 ;
        RECT 64.945 105.455 66.255 105.755 ;
        RECT 65.680 105.420 66.060 105.455 ;
        RECT 82.775 105.440 83.865 105.820 ;
        RECT 87.260 105.445 100.110 105.780 ;
        RECT 104.275 105.775 104.655 105.820 ;
        RECT 103.540 105.475 104.850 105.775 ;
        RECT 123.645 105.490 127.795 105.760 ;
        RECT 104.275 105.440 104.655 105.475 ;
        RECT 73.335 104.910 106.285 104.945 ;
        RECT 41.035 104.580 106.285 104.910 ;
        RECT 41.035 104.560 74.115 104.580 ;
        RECT 108.080 104.570 112.340 104.925 ;
        RECT 40.905 97.370 78.455 97.395 ;
        RECT 40.905 97.110 106.530 97.370 ;
        RECT 77.755 97.085 106.530 97.110 ;
        RECT 108.200 97.065 114.905 97.365 ;
        RECT 44.610 96.200 45.810 96.580 ;
        RECT 64.135 96.300 65.370 96.680 ;
        RECT 81.060 96.175 82.515 96.555 ;
        RECT 104.755 96.275 106.035 96.655 ;
        RECT 65.550 95.945 65.930 95.980 ;
        RECT 44.050 95.840 44.430 95.880 ;
        RECT 43.980 95.535 46.815 95.840 ;
        RECT 62.795 95.635 65.930 95.945 ;
        RECT 104.195 95.920 104.575 95.955 ;
        RECT 82.695 95.815 83.075 95.855 ;
        RECT 65.550 95.600 65.930 95.635 ;
        RECT 44.050 95.500 44.430 95.535 ;
        RECT 82.625 95.510 85.460 95.815 ;
        RECT 101.440 95.610 104.575 95.920 ;
        RECT 123.705 95.895 130.445 96.195 ;
        RECT 104.195 95.575 104.575 95.610 ;
        RECT 82.695 95.475 83.075 95.510 ;
        RECT 14.380 93.925 14.760 94.305 ;
        RECT 21.280 93.915 21.660 94.295 ;
        RECT 26.095 94.125 29.500 94.565 ;
        RECT 29.840 93.925 30.220 94.305 ;
        RECT 32.555 93.965 32.935 94.345 ;
        RECT 36.740 93.915 37.120 94.295 ;
        RECT 44.610 93.900 47.870 94.280 ;
        RECT 48.610 93.900 51.870 94.280 ;
        RECT 58.110 93.900 61.370 94.280 ;
        RECT 62.110 93.900 65.370 94.280 ;
        RECT 11.705 93.500 13.445 93.790 ;
        RECT 18.205 93.420 20.815 93.845 ;
        RECT 27.165 93.500 28.905 93.790 ;
        RECT 30.955 93.450 32.155 93.740 ;
        RECT 33.665 93.420 36.260 93.795 ;
        RECT 37.875 93.515 38.255 93.895 ;
        RECT 81.220 93.875 82.515 94.255 ;
        RECT 87.255 93.875 90.515 94.255 ;
        RECT 91.255 93.875 92.440 94.255 ;
        RECT 94.705 93.875 96.015 94.255 ;
        RECT 96.755 93.875 100.015 94.255 ;
        RECT 104.755 93.875 105.770 94.255 ;
        RECT 108.835 94.120 112.250 94.540 ;
        RECT 112.580 93.900 112.960 94.280 ;
        RECT 115.295 93.940 115.675 94.320 ;
        RECT 119.480 93.890 119.860 94.270 ;
        RECT 124.295 94.100 127.750 94.540 ;
        RECT 130.755 93.940 131.135 94.320 ;
        RECT 44.050 93.200 44.430 93.580 ;
        RECT 48.050 93.200 48.430 93.580 ;
        RECT 52.050 93.535 52.430 93.580 ;
        RECT 57.550 93.535 57.930 93.580 ;
        RECT 52.000 93.220 57.935 93.535 ;
        RECT 52.050 93.200 52.430 93.220 ;
        RECT 57.550 93.200 57.930 93.220 ;
        RECT 61.550 93.200 61.930 93.580 ;
        RECT 65.550 93.200 65.930 93.580 ;
        RECT 82.695 93.175 83.075 93.555 ;
        RECT 86.695 93.175 87.075 93.555 ;
        RECT 90.695 93.510 91.075 93.555 ;
        RECT 96.195 93.510 96.575 93.555 ;
        RECT 90.645 93.195 96.580 93.510 ;
        RECT 90.695 93.175 91.075 93.195 ;
        RECT 96.195 93.175 96.575 93.195 ;
        RECT 100.195 93.175 100.575 93.555 ;
        RECT 104.195 93.175 104.575 93.555 ;
        RECT 109.905 93.475 111.645 93.765 ;
        RECT 113.695 93.425 114.895 93.715 ;
        RECT 116.405 93.385 119.035 93.840 ;
        RECT 120.615 93.490 120.995 93.870 ;
        RECT 129.155 93.425 130.355 93.715 ;
        RECT 136.075 93.490 136.455 93.870 ;
        RECT 74.785 92.550 95.560 92.925 ;
        RECT 123.110 92.715 139.030 93.015 ;
        RECT 45.275 91.985 72.585 92.325 ;
        RECT 123.645 91.970 140.590 92.270 ;
        RECT 24.890 91.280 32.150 91.580 ;
        RECT 20.390 90.980 23.495 91.255 ;
        RECT 25.445 90.745 29.530 91.015 ;
        RECT 35.850 90.980 39.600 91.255 ;
        RECT 73.815 91.195 105.780 91.585 ;
        RECT 118.590 90.955 121.720 91.230 ;
        RECT 40.905 90.855 59.575 90.865 ;
        RECT 40.905 90.840 70.925 90.855 ;
        RECT 40.905 90.830 98.220 90.840 ;
        RECT 40.905 90.545 107.225 90.830 ;
        RECT 70.660 90.520 107.225 90.545 ;
        RECT 124.840 90.060 128.970 90.360 ;
        RECT 131.345 90.010 135.845 90.320 ;
        RECT 40.375 89.850 76.285 89.875 ;
        RECT 29.105 89.485 35.495 89.775 ;
        RECT 40.375 89.605 107.625 89.850 ;
        RECT 75.880 89.580 107.625 89.605 ;
        RECT 111.845 89.460 118.235 89.750 ;
        RECT 127.305 89.460 133.695 89.750 ;
        RECT 13.060 88.905 23.715 89.240 ;
        RECT 28.520 88.905 39.025 89.240 ;
        RECT 63.995 89.040 74.545 89.375 ;
        RECT 111.260 88.880 121.740 89.215 ;
        RECT 44.590 88.400 47.890 88.780 ;
        RECT 48.590 88.400 51.890 88.780 ;
        RECT 58.090 88.400 61.390 88.780 ;
        RECT 62.090 88.400 65.390 88.780 ;
        RECT 81.230 88.375 82.535 88.755 ;
        RECT 87.235 88.375 90.535 88.755 ;
        RECT 91.235 88.375 92.595 88.755 ;
        RECT 94.570 88.375 96.035 88.755 ;
        RECT 96.735 88.375 100.035 88.755 ;
        RECT 104.735 88.375 105.915 88.755 ;
        RECT 126.070 88.295 128.990 88.595 ;
        RECT 132.535 88.280 135.905 88.580 ;
        RECT 44.050 88.055 44.430 88.090 ;
        RECT 13.030 87.585 14.810 87.875 ;
        RECT 20.405 87.555 21.715 87.875 ;
        RECT 26.085 87.570 26.465 87.950 ;
        RECT 28.490 87.585 30.270 87.875 ;
        RECT 31.745 87.675 32.935 87.960 ;
        RECT 35.865 87.555 37.175 87.875 ;
        RECT 43.785 87.745 46.795 88.055 ;
        RECT 44.050 87.710 44.430 87.745 ;
        RECT 48.050 87.710 49.140 88.090 ;
        RECT 52.050 88.085 52.430 88.090 ;
        RECT 49.570 87.720 52.435 88.085 ;
        RECT 57.550 88.065 57.930 88.090 ;
        RECT 57.535 87.745 59.680 88.065 ;
        RECT 52.050 87.710 52.430 87.720 ;
        RECT 57.550 87.710 57.930 87.745 ;
        RECT 60.595 87.710 61.930 88.090 ;
        RECT 65.550 88.070 65.930 88.090 ;
        RECT 63.085 87.750 65.995 88.070 ;
        RECT 82.695 88.030 83.075 88.065 ;
        RECT 65.550 87.710 65.930 87.750 ;
        RECT 82.430 87.720 85.440 88.030 ;
        RECT 82.695 87.685 83.075 87.720 ;
        RECT 86.695 87.685 87.785 88.065 ;
        RECT 90.695 88.060 91.075 88.065 ;
        RECT 88.215 87.695 91.080 88.060 ;
        RECT 96.195 88.040 96.575 88.065 ;
        RECT 96.180 87.720 98.325 88.040 ;
        RECT 90.695 87.685 91.075 87.695 ;
        RECT 96.195 87.685 96.575 87.720 ;
        RECT 99.240 87.685 100.575 88.065 ;
        RECT 104.195 88.045 104.575 88.065 ;
        RECT 101.730 87.725 104.640 88.045 ;
        RECT 104.195 87.685 104.575 87.725 ;
        RECT 108.825 87.545 109.205 87.925 ;
        RECT 111.230 87.560 113.010 87.850 ;
        RECT 114.485 87.650 115.675 87.935 ;
        RECT 118.605 87.530 119.915 87.850 ;
        RECT 124.285 87.545 124.665 87.925 ;
        RECT 129.945 87.650 131.135 87.935 ;
        RECT 11.760 86.970 12.140 87.350 ;
        RECT 18.215 87.000 18.595 87.380 ;
        RECT 27.220 86.970 27.600 87.350 ;
        RECT 30.965 87.010 31.345 87.390 ;
        RECT 33.675 87.000 34.055 87.380 ;
        RECT 35.085 86.845 38.265 87.165 ;
        RECT 109.960 86.945 110.340 87.325 ;
        RECT 113.705 86.985 114.085 87.365 ;
        RECT 116.415 86.975 116.795 87.355 ;
        RECT 117.825 86.820 121.005 87.140 ;
        RECT 129.165 86.985 129.545 87.365 ;
        RECT 133.285 86.820 136.465 87.140 ;
        RECT 44.590 86.400 45.875 86.780 ;
        RECT 63.905 86.400 65.390 86.780 ;
        RECT 81.045 86.375 82.535 86.755 ;
        RECT 104.735 86.375 105.810 86.755 ;
        RECT 44.050 85.710 45.140 86.090 ;
        RECT 48.535 85.715 61.385 86.050 ;
        RECT 65.550 86.045 65.930 86.090 ;
        RECT 64.815 85.745 66.125 86.045 ;
        RECT 65.550 85.710 65.930 85.745 ;
        RECT 82.695 85.685 83.785 86.065 ;
        RECT 87.180 85.690 100.030 86.025 ;
        RECT 104.195 86.020 104.575 86.065 ;
        RECT 103.460 85.720 104.770 86.020 ;
        RECT 123.565 85.735 127.715 86.005 ;
        RECT 104.195 85.685 104.575 85.720 ;
        RECT 40.905 85.190 73.985 85.200 ;
        RECT 40.905 84.850 106.205 85.190 ;
        RECT 73.255 84.825 106.205 84.850 ;
        RECT 108.000 84.815 112.260 85.170 ;
        RECT 77.860 77.635 106.635 77.655 ;
        RECT 41.035 77.370 106.635 77.635 ;
        RECT 41.035 77.350 78.585 77.370 ;
        RECT 108.305 77.350 115.010 77.650 ;
        RECT 44.740 76.440 45.940 76.820 ;
        RECT 64.265 76.540 65.500 76.920 ;
        RECT 81.165 76.460 82.620 76.840 ;
        RECT 104.860 76.560 106.140 76.940 ;
        RECT 65.680 76.185 66.060 76.220 ;
        RECT 104.300 76.205 104.680 76.240 ;
        RECT 44.180 76.080 44.560 76.120 ;
        RECT 44.110 75.775 46.945 76.080 ;
        RECT 62.925 75.875 66.060 76.185 ;
        RECT 82.800 76.100 83.180 76.140 ;
        RECT 65.680 75.840 66.060 75.875 ;
        RECT 82.730 75.795 85.565 76.100 ;
        RECT 101.545 75.895 104.680 76.205 ;
        RECT 123.810 76.180 130.550 76.480 ;
        RECT 104.300 75.860 104.680 75.895 ;
        RECT 44.180 75.740 44.560 75.775 ;
        RECT 82.800 75.760 83.180 75.795 ;
        RECT 14.510 74.165 14.890 74.545 ;
        RECT 21.410 74.155 21.790 74.535 ;
        RECT 26.225 74.365 29.630 74.805 ;
        RECT 29.970 74.165 30.350 74.545 ;
        RECT 32.685 74.205 33.065 74.585 ;
        RECT 36.870 74.155 37.250 74.535 ;
        RECT 44.740 74.140 48.000 74.520 ;
        RECT 48.740 74.140 52.000 74.520 ;
        RECT 58.240 74.140 61.500 74.520 ;
        RECT 62.240 74.140 65.500 74.520 ;
        RECT 81.325 74.160 82.620 74.540 ;
        RECT 87.360 74.160 90.620 74.540 ;
        RECT 91.360 74.160 92.545 74.540 ;
        RECT 94.810 74.160 96.120 74.540 ;
        RECT 96.860 74.160 100.120 74.540 ;
        RECT 104.860 74.160 105.875 74.540 ;
        RECT 108.940 74.405 112.355 74.825 ;
        RECT 112.685 74.185 113.065 74.565 ;
        RECT 115.400 74.225 115.780 74.605 ;
        RECT 119.585 74.175 119.965 74.555 ;
        RECT 124.400 74.385 127.855 74.825 ;
        RECT 130.860 74.225 131.240 74.605 ;
        RECT 11.835 73.740 13.575 74.030 ;
        RECT 18.335 73.660 20.945 74.085 ;
        RECT 27.295 73.740 29.035 74.030 ;
        RECT 31.085 73.690 32.285 73.980 ;
        RECT 33.795 73.660 36.390 74.035 ;
        RECT 38.005 73.755 38.385 74.135 ;
        RECT 44.180 73.440 44.560 73.820 ;
        RECT 48.180 73.440 48.560 73.820 ;
        RECT 52.180 73.775 52.560 73.820 ;
        RECT 57.680 73.775 58.060 73.820 ;
        RECT 52.130 73.460 58.065 73.775 ;
        RECT 52.180 73.440 52.560 73.460 ;
        RECT 57.680 73.440 58.060 73.460 ;
        RECT 61.680 73.440 62.060 73.820 ;
        RECT 65.680 73.440 66.060 73.820 ;
        RECT 82.800 73.460 83.180 73.840 ;
        RECT 86.800 73.460 87.180 73.840 ;
        RECT 90.800 73.795 91.180 73.840 ;
        RECT 96.300 73.795 96.680 73.840 ;
        RECT 90.750 73.480 96.685 73.795 ;
        RECT 90.800 73.460 91.180 73.480 ;
        RECT 96.300 73.460 96.680 73.480 ;
        RECT 100.300 73.460 100.680 73.840 ;
        RECT 104.300 73.460 104.680 73.840 ;
        RECT 110.010 73.760 111.750 74.050 ;
        RECT 113.800 73.710 115.000 74.000 ;
        RECT 116.510 73.670 119.140 74.125 ;
        RECT 120.720 73.775 121.100 74.155 ;
        RECT 129.260 73.710 130.460 74.000 ;
        RECT 136.180 73.775 136.560 74.155 ;
        RECT 74.890 72.835 95.665 73.210 ;
        RECT 123.215 73.000 139.135 73.300 ;
        RECT 45.405 72.225 72.715 72.565 ;
        RECT 123.750 72.255 140.695 72.555 ;
        RECT 25.020 71.520 32.280 71.820 ;
        RECT 20.520 71.220 23.625 71.495 ;
        RECT 25.575 70.985 29.660 71.255 ;
        RECT 35.980 71.220 39.730 71.495 ;
        RECT 73.920 71.480 105.885 71.870 ;
        RECT 118.695 71.240 121.825 71.515 ;
        RECT 70.765 71.115 98.325 71.125 ;
        RECT 41.035 71.095 59.705 71.105 ;
        RECT 70.765 71.095 107.330 71.115 ;
        RECT 41.035 70.805 107.330 71.095 ;
        RECT 41.035 70.785 71.055 70.805 ;
        RECT 124.945 70.345 129.075 70.645 ;
        RECT 131.450 70.295 135.950 70.605 ;
        RECT 75.985 70.115 107.730 70.135 ;
        RECT 29.235 69.725 35.625 70.015 ;
        RECT 40.505 69.865 107.730 70.115 ;
        RECT 40.505 69.845 76.415 69.865 ;
        RECT 111.950 69.745 118.340 70.035 ;
        RECT 127.410 69.745 133.800 70.035 ;
        RECT 13.190 69.145 23.845 69.480 ;
        RECT 28.650 69.145 39.155 69.480 ;
        RECT 64.125 69.280 74.675 69.615 ;
        RECT 111.365 69.165 121.845 69.500 ;
        RECT 44.720 68.640 48.020 69.020 ;
        RECT 48.720 68.640 52.020 69.020 ;
        RECT 58.220 68.640 61.520 69.020 ;
        RECT 62.220 68.640 65.520 69.020 ;
        RECT 81.335 68.660 82.640 69.040 ;
        RECT 87.340 68.660 90.640 69.040 ;
        RECT 91.340 68.660 92.700 69.040 ;
        RECT 94.675 68.660 96.140 69.040 ;
        RECT 96.840 68.660 100.140 69.040 ;
        RECT 104.840 68.660 106.020 69.040 ;
        RECT 126.175 68.580 129.095 68.880 ;
        RECT 132.640 68.565 136.010 68.865 ;
        RECT 44.180 68.295 44.560 68.330 ;
        RECT 13.160 67.825 14.940 68.115 ;
        RECT 20.535 67.795 21.845 68.115 ;
        RECT 26.215 67.810 26.595 68.190 ;
        RECT 28.620 67.825 30.400 68.115 ;
        RECT 31.875 67.915 33.065 68.200 ;
        RECT 35.995 67.795 37.305 68.115 ;
        RECT 43.915 67.985 46.925 68.295 ;
        RECT 44.180 67.950 44.560 67.985 ;
        RECT 48.180 67.950 49.270 68.330 ;
        RECT 52.180 68.325 52.560 68.330 ;
        RECT 49.700 67.960 52.565 68.325 ;
        RECT 57.680 68.305 58.060 68.330 ;
        RECT 57.665 67.985 59.810 68.305 ;
        RECT 52.180 67.950 52.560 67.960 ;
        RECT 57.680 67.950 58.060 67.985 ;
        RECT 60.725 67.950 62.060 68.330 ;
        RECT 65.680 68.310 66.060 68.330 ;
        RECT 82.800 68.315 83.180 68.350 ;
        RECT 63.215 67.990 66.125 68.310 ;
        RECT 82.535 68.005 85.545 68.315 ;
        RECT 65.680 67.950 66.060 67.990 ;
        RECT 82.800 67.970 83.180 68.005 ;
        RECT 86.800 67.970 87.890 68.350 ;
        RECT 90.800 68.345 91.180 68.350 ;
        RECT 88.320 67.980 91.185 68.345 ;
        RECT 96.300 68.325 96.680 68.350 ;
        RECT 96.285 68.005 98.430 68.325 ;
        RECT 90.800 67.970 91.180 67.980 ;
        RECT 96.300 67.970 96.680 68.005 ;
        RECT 99.345 67.970 100.680 68.350 ;
        RECT 104.300 68.330 104.680 68.350 ;
        RECT 101.835 68.010 104.745 68.330 ;
        RECT 104.300 67.970 104.680 68.010 ;
        RECT 108.930 67.830 109.310 68.210 ;
        RECT 111.335 67.845 113.115 68.135 ;
        RECT 114.590 67.935 115.780 68.220 ;
        RECT 118.710 67.815 120.020 68.135 ;
        RECT 124.390 67.830 124.770 68.210 ;
        RECT 130.050 67.935 131.240 68.220 ;
        RECT 11.890 67.210 12.270 67.590 ;
        RECT 18.345 67.240 18.725 67.620 ;
        RECT 27.350 67.210 27.730 67.590 ;
        RECT 31.095 67.250 31.475 67.630 ;
        RECT 33.805 67.240 34.185 67.620 ;
        RECT 35.215 67.085 38.395 67.405 ;
        RECT 110.065 67.230 110.445 67.610 ;
        RECT 113.810 67.270 114.190 67.650 ;
        RECT 116.520 67.260 116.900 67.640 ;
        RECT 117.930 67.105 121.110 67.425 ;
        RECT 129.270 67.270 129.650 67.650 ;
        RECT 133.390 67.105 136.570 67.425 ;
        RECT 44.720 66.640 46.005 67.020 ;
        RECT 64.035 66.640 65.520 67.020 ;
        RECT 81.150 66.660 82.640 67.040 ;
        RECT 104.840 66.660 105.915 67.040 ;
        RECT 44.180 65.950 45.270 66.330 ;
        RECT 48.665 65.955 61.515 66.290 ;
        RECT 65.680 66.285 66.060 66.330 ;
        RECT 64.945 65.985 66.255 66.285 ;
        RECT 65.680 65.950 66.060 65.985 ;
        RECT 82.800 65.970 83.890 66.350 ;
        RECT 87.285 65.975 100.135 66.310 ;
        RECT 104.300 66.305 104.680 66.350 ;
        RECT 103.565 66.005 104.875 66.305 ;
        RECT 123.670 66.020 127.820 66.290 ;
        RECT 104.300 65.970 104.680 66.005 ;
        RECT 73.360 65.440 106.310 65.475 ;
        RECT 41.035 65.110 106.310 65.440 ;
        RECT 41.035 65.090 74.115 65.110 ;
        RECT 108.105 65.100 112.365 65.455 ;
        RECT 40.985 57.685 78.535 57.825 ;
        RECT 40.985 57.540 106.635 57.685 ;
        RECT 77.860 57.400 106.635 57.540 ;
        RECT 108.305 57.380 115.010 57.680 ;
        RECT 44.690 56.630 45.890 57.010 ;
        RECT 64.215 56.730 65.450 57.110 ;
        RECT 81.165 56.490 82.620 56.870 ;
        RECT 104.860 56.590 106.140 56.970 ;
        RECT 65.630 56.375 66.010 56.410 ;
        RECT 44.130 56.270 44.510 56.310 ;
        RECT 44.060 55.965 46.895 56.270 ;
        RECT 62.875 56.065 66.010 56.375 ;
        RECT 104.300 56.235 104.680 56.270 ;
        RECT 82.800 56.130 83.180 56.170 ;
        RECT 65.630 56.030 66.010 56.065 ;
        RECT 44.130 55.930 44.510 55.965 ;
        RECT 82.730 55.825 85.565 56.130 ;
        RECT 101.545 55.925 104.680 56.235 ;
        RECT 123.810 56.210 130.550 56.510 ;
        RECT 104.300 55.890 104.680 55.925 ;
        RECT 82.800 55.790 83.180 55.825 ;
        RECT 14.460 54.355 14.840 54.735 ;
        RECT 21.360 54.345 21.740 54.725 ;
        RECT 26.175 54.555 29.580 54.995 ;
        RECT 29.920 54.355 30.300 54.735 ;
        RECT 32.635 54.395 33.015 54.775 ;
        RECT 36.820 54.345 37.200 54.725 ;
        RECT 44.690 54.330 47.950 54.710 ;
        RECT 48.690 54.330 51.950 54.710 ;
        RECT 58.190 54.330 61.450 54.710 ;
        RECT 62.190 54.330 65.450 54.710 ;
        RECT 11.785 53.930 13.525 54.220 ;
        RECT 18.285 53.850 20.895 54.275 ;
        RECT 27.245 53.930 28.985 54.220 ;
        RECT 31.035 53.880 32.235 54.170 ;
        RECT 33.745 53.850 36.340 54.225 ;
        RECT 37.955 53.945 38.335 54.325 ;
        RECT 81.325 54.190 82.620 54.570 ;
        RECT 87.360 54.190 90.620 54.570 ;
        RECT 91.360 54.190 92.545 54.570 ;
        RECT 94.810 54.190 96.120 54.570 ;
        RECT 96.860 54.190 100.120 54.570 ;
        RECT 104.860 54.190 105.875 54.570 ;
        RECT 108.940 54.435 112.355 54.855 ;
        RECT 112.685 54.215 113.065 54.595 ;
        RECT 115.400 54.255 115.780 54.635 ;
        RECT 119.585 54.205 119.965 54.585 ;
        RECT 124.400 54.415 127.855 54.855 ;
        RECT 130.860 54.255 131.240 54.635 ;
        RECT 44.130 53.630 44.510 54.010 ;
        RECT 48.130 53.630 48.510 54.010 ;
        RECT 52.130 53.965 52.510 54.010 ;
        RECT 57.630 53.965 58.010 54.010 ;
        RECT 52.080 53.650 58.015 53.965 ;
        RECT 52.130 53.630 52.510 53.650 ;
        RECT 57.630 53.630 58.010 53.650 ;
        RECT 61.630 53.630 62.010 54.010 ;
        RECT 65.630 53.630 66.010 54.010 ;
        RECT 82.800 53.490 83.180 53.870 ;
        RECT 86.800 53.490 87.180 53.870 ;
        RECT 90.800 53.825 91.180 53.870 ;
        RECT 96.300 53.825 96.680 53.870 ;
        RECT 90.750 53.510 96.685 53.825 ;
        RECT 90.800 53.490 91.180 53.510 ;
        RECT 96.300 53.490 96.680 53.510 ;
        RECT 100.300 53.490 100.680 53.870 ;
        RECT 104.300 53.490 104.680 53.870 ;
        RECT 110.010 53.790 111.750 54.080 ;
        RECT 113.800 53.740 115.000 54.030 ;
        RECT 116.510 53.700 119.140 54.155 ;
        RECT 120.720 53.805 121.100 54.185 ;
        RECT 129.260 53.740 130.460 54.030 ;
        RECT 136.180 53.805 136.560 54.185 ;
        RECT 74.890 52.865 95.665 53.240 ;
        RECT 123.215 53.030 139.135 53.330 ;
        RECT 45.355 52.415 72.665 52.755 ;
        RECT 123.750 52.285 140.695 52.585 ;
        RECT 24.970 51.710 32.230 52.010 ;
        RECT 20.470 51.410 23.575 51.685 ;
        RECT 25.525 51.175 29.610 51.445 ;
        RECT 35.930 51.410 39.680 51.685 ;
        RECT 73.920 51.510 105.885 51.900 ;
        RECT 40.985 51.285 59.655 51.295 ;
        RECT 40.985 51.155 71.005 51.285 ;
        RECT 118.695 51.270 121.825 51.545 ;
        RECT 40.985 51.145 98.325 51.155 ;
        RECT 40.985 50.975 107.330 51.145 ;
        RECT 70.765 50.835 107.330 50.975 ;
        RECT 124.945 50.375 129.075 50.675 ;
        RECT 131.450 50.325 135.950 50.635 ;
        RECT 29.185 49.915 35.575 50.205 ;
        RECT 40.455 50.165 76.365 50.305 ;
        RECT 40.455 50.035 107.730 50.165 ;
        RECT 75.985 49.895 107.730 50.035 ;
        RECT 13.140 49.335 23.795 49.670 ;
        RECT 28.600 49.335 39.105 49.670 ;
        RECT 64.075 49.470 74.625 49.805 ;
        RECT 111.950 49.775 118.340 50.065 ;
        RECT 127.410 49.775 133.800 50.065 ;
        RECT 44.670 48.830 47.970 49.210 ;
        RECT 48.670 48.830 51.970 49.210 ;
        RECT 58.170 48.830 61.470 49.210 ;
        RECT 62.170 48.830 65.470 49.210 ;
        RECT 111.365 49.195 121.845 49.530 ;
        RECT 81.335 48.690 82.640 49.070 ;
        RECT 87.340 48.690 90.640 49.070 ;
        RECT 91.340 48.690 92.700 49.070 ;
        RECT 94.675 48.690 96.140 49.070 ;
        RECT 96.840 48.690 100.140 49.070 ;
        RECT 104.840 48.690 106.020 49.070 ;
        RECT 126.175 48.610 129.095 48.910 ;
        RECT 132.640 48.595 136.010 48.895 ;
        RECT 44.130 48.485 44.510 48.520 ;
        RECT 13.110 48.015 14.890 48.305 ;
        RECT 20.485 47.985 21.795 48.305 ;
        RECT 26.165 48.000 26.545 48.380 ;
        RECT 28.570 48.015 30.350 48.305 ;
        RECT 31.825 48.105 33.015 48.390 ;
        RECT 35.945 47.985 37.255 48.305 ;
        RECT 43.865 48.175 46.875 48.485 ;
        RECT 44.130 48.140 44.510 48.175 ;
        RECT 48.130 48.140 49.220 48.520 ;
        RECT 52.130 48.515 52.510 48.520 ;
        RECT 49.650 48.150 52.515 48.515 ;
        RECT 57.630 48.495 58.010 48.520 ;
        RECT 57.615 48.175 59.760 48.495 ;
        RECT 52.130 48.140 52.510 48.150 ;
        RECT 57.630 48.140 58.010 48.175 ;
        RECT 60.675 48.140 62.010 48.520 ;
        RECT 65.630 48.500 66.010 48.520 ;
        RECT 63.165 48.180 66.075 48.500 ;
        RECT 82.800 48.345 83.180 48.380 ;
        RECT 65.630 48.140 66.010 48.180 ;
        RECT 82.535 48.035 85.545 48.345 ;
        RECT 82.800 48.000 83.180 48.035 ;
        RECT 86.800 48.000 87.890 48.380 ;
        RECT 90.800 48.375 91.180 48.380 ;
        RECT 88.320 48.010 91.185 48.375 ;
        RECT 96.300 48.355 96.680 48.380 ;
        RECT 96.285 48.035 98.430 48.355 ;
        RECT 90.800 48.000 91.180 48.010 ;
        RECT 96.300 48.000 96.680 48.035 ;
        RECT 99.345 48.000 100.680 48.380 ;
        RECT 104.300 48.360 104.680 48.380 ;
        RECT 101.835 48.040 104.745 48.360 ;
        RECT 104.300 48.000 104.680 48.040 ;
        RECT 108.930 47.860 109.310 48.240 ;
        RECT 111.335 47.875 113.115 48.165 ;
        RECT 114.590 47.965 115.780 48.250 ;
        RECT 118.710 47.845 120.020 48.165 ;
        RECT 124.390 47.860 124.770 48.240 ;
        RECT 130.050 47.965 131.240 48.250 ;
        RECT 11.840 47.400 12.220 47.780 ;
        RECT 18.295 47.430 18.675 47.810 ;
        RECT 27.300 47.400 27.680 47.780 ;
        RECT 31.045 47.440 31.425 47.820 ;
        RECT 33.755 47.430 34.135 47.810 ;
        RECT 35.165 47.275 38.345 47.595 ;
        RECT 110.065 47.260 110.445 47.640 ;
        RECT 113.810 47.300 114.190 47.680 ;
        RECT 116.520 47.290 116.900 47.670 ;
        RECT 44.670 46.830 45.955 47.210 ;
        RECT 63.985 46.830 65.470 47.210 ;
        RECT 117.930 47.135 121.110 47.455 ;
        RECT 129.270 47.300 129.650 47.680 ;
        RECT 133.390 47.135 136.570 47.455 ;
        RECT 81.150 46.690 82.640 47.070 ;
        RECT 104.840 46.690 105.915 47.070 ;
        RECT 44.130 46.140 45.220 46.520 ;
        RECT 48.615 46.145 61.465 46.480 ;
        RECT 65.630 46.475 66.010 46.520 ;
        RECT 64.895 46.175 66.205 46.475 ;
        RECT 65.630 46.140 66.010 46.175 ;
        RECT 82.800 46.000 83.890 46.380 ;
        RECT 87.285 46.005 100.135 46.340 ;
        RECT 104.300 46.335 104.680 46.380 ;
        RECT 103.565 46.035 104.875 46.335 ;
        RECT 123.670 46.050 127.820 46.320 ;
        RECT 104.300 46.000 104.680 46.035 ;
        RECT 40.985 45.505 74.065 45.630 ;
        RECT 40.985 45.280 106.310 45.505 ;
        RECT 73.360 45.140 106.310 45.280 ;
        RECT 108.105 45.130 112.365 45.485 ;
        RECT 40.955 38.020 78.505 38.030 ;
        RECT 40.955 37.745 106.635 38.020 ;
        RECT 77.860 37.735 106.635 37.745 ;
        RECT 108.305 37.715 115.010 38.015 ;
        RECT 44.660 36.835 45.860 37.215 ;
        RECT 64.185 36.935 65.420 37.315 ;
        RECT 81.165 36.825 82.620 37.205 ;
        RECT 104.860 36.925 106.140 37.305 ;
        RECT 65.600 36.580 65.980 36.615 ;
        RECT 44.100 36.475 44.480 36.515 ;
        RECT 44.030 36.170 46.865 36.475 ;
        RECT 62.845 36.270 65.980 36.580 ;
        RECT 104.300 36.570 104.680 36.605 ;
        RECT 82.800 36.465 83.180 36.505 ;
        RECT 65.600 36.235 65.980 36.270 ;
        RECT 44.100 36.135 44.480 36.170 ;
        RECT 82.730 36.160 85.565 36.465 ;
        RECT 101.545 36.260 104.680 36.570 ;
        RECT 123.810 36.545 130.550 36.845 ;
        RECT 104.300 36.225 104.680 36.260 ;
        RECT 82.800 36.125 83.180 36.160 ;
        RECT 14.430 34.560 14.810 34.940 ;
        RECT 21.330 34.550 21.710 34.930 ;
        RECT 26.145 34.760 29.550 35.200 ;
        RECT 29.890 34.560 30.270 34.940 ;
        RECT 32.605 34.600 32.985 34.980 ;
        RECT 36.790 34.550 37.170 34.930 ;
        RECT 44.660 34.535 47.920 34.915 ;
        RECT 48.660 34.535 51.920 34.915 ;
        RECT 58.160 34.535 61.420 34.915 ;
        RECT 62.160 34.535 65.420 34.915 ;
        RECT 11.755 34.135 13.495 34.425 ;
        RECT 18.255 34.055 20.865 34.480 ;
        RECT 27.215 34.135 28.955 34.425 ;
        RECT 31.005 34.085 32.205 34.375 ;
        RECT 33.715 34.055 36.310 34.430 ;
        RECT 37.925 34.150 38.305 34.530 ;
        RECT 81.325 34.525 82.620 34.905 ;
        RECT 87.360 34.525 90.620 34.905 ;
        RECT 91.360 34.525 92.545 34.905 ;
        RECT 94.810 34.525 96.120 34.905 ;
        RECT 96.860 34.525 100.120 34.905 ;
        RECT 104.860 34.525 105.875 34.905 ;
        RECT 108.940 34.770 112.355 35.190 ;
        RECT 112.685 34.550 113.065 34.930 ;
        RECT 115.400 34.590 115.780 34.970 ;
        RECT 119.585 34.540 119.965 34.920 ;
        RECT 124.400 34.750 127.855 35.190 ;
        RECT 130.860 34.590 131.240 34.970 ;
        RECT 44.100 33.835 44.480 34.215 ;
        RECT 48.100 33.835 48.480 34.215 ;
        RECT 52.100 34.170 52.480 34.215 ;
        RECT 57.600 34.170 57.980 34.215 ;
        RECT 52.050 33.855 57.985 34.170 ;
        RECT 52.100 33.835 52.480 33.855 ;
        RECT 57.600 33.835 57.980 33.855 ;
        RECT 61.600 33.835 61.980 34.215 ;
        RECT 65.600 33.835 65.980 34.215 ;
        RECT 82.800 33.825 83.180 34.205 ;
        RECT 86.800 33.825 87.180 34.205 ;
        RECT 90.800 34.160 91.180 34.205 ;
        RECT 96.300 34.160 96.680 34.205 ;
        RECT 90.750 33.845 96.685 34.160 ;
        RECT 90.800 33.825 91.180 33.845 ;
        RECT 96.300 33.825 96.680 33.845 ;
        RECT 100.300 33.825 100.680 34.205 ;
        RECT 104.300 33.825 104.680 34.205 ;
        RECT 110.010 34.125 111.750 34.415 ;
        RECT 113.800 34.075 115.000 34.365 ;
        RECT 116.510 34.035 119.140 34.490 ;
        RECT 120.720 34.140 121.100 34.520 ;
        RECT 129.260 34.075 130.460 34.365 ;
        RECT 136.180 34.140 136.560 34.520 ;
        RECT 74.890 33.200 95.665 33.575 ;
        RECT 123.215 33.365 139.135 33.665 ;
        RECT 45.325 32.620 72.635 32.960 ;
        RECT 123.750 32.620 140.695 32.920 ;
        RECT 24.940 31.915 32.200 32.215 ;
        RECT 20.440 31.615 23.545 31.890 ;
        RECT 25.495 31.380 29.580 31.650 ;
        RECT 35.900 31.615 39.650 31.890 ;
        RECT 73.920 31.845 105.885 32.235 ;
        RECT 118.695 31.605 121.825 31.880 ;
        RECT 40.955 31.490 59.625 31.500 ;
        RECT 40.955 31.480 98.325 31.490 ;
        RECT 40.955 31.180 107.330 31.480 ;
        RECT 70.765 31.170 107.330 31.180 ;
        RECT 124.945 30.710 129.075 31.010 ;
        RECT 131.450 30.660 135.950 30.970 ;
        RECT 40.425 30.500 76.335 30.510 ;
        RECT 29.155 30.120 35.545 30.410 ;
        RECT 40.425 30.240 107.730 30.500 ;
        RECT 75.985 30.230 107.730 30.240 ;
        RECT 111.950 30.110 118.340 30.400 ;
        RECT 127.410 30.110 133.800 30.400 ;
        RECT 13.110 29.540 23.765 29.875 ;
        RECT 28.570 29.540 39.075 29.875 ;
        RECT 64.045 29.675 74.595 30.010 ;
        RECT 111.365 29.530 121.845 29.865 ;
        RECT 44.640 29.035 47.940 29.415 ;
        RECT 48.640 29.035 51.940 29.415 ;
        RECT 58.140 29.035 61.440 29.415 ;
        RECT 62.140 29.035 65.440 29.415 ;
        RECT 81.335 29.025 82.640 29.405 ;
        RECT 87.340 29.025 90.640 29.405 ;
        RECT 91.340 29.025 92.700 29.405 ;
        RECT 94.675 29.025 96.140 29.405 ;
        RECT 96.840 29.025 100.140 29.405 ;
        RECT 104.840 29.025 106.020 29.405 ;
        RECT 126.175 28.945 129.095 29.245 ;
        RECT 132.640 28.930 136.010 29.230 ;
        RECT 44.100 28.690 44.480 28.725 ;
        RECT 13.080 28.220 14.860 28.510 ;
        RECT 20.455 28.190 21.765 28.510 ;
        RECT 26.135 28.205 26.515 28.585 ;
        RECT 28.540 28.220 30.320 28.510 ;
        RECT 31.795 28.310 32.985 28.595 ;
        RECT 35.915 28.190 37.225 28.510 ;
        RECT 43.835 28.380 46.845 28.690 ;
        RECT 44.100 28.345 44.480 28.380 ;
        RECT 48.100 28.345 49.190 28.725 ;
        RECT 52.100 28.720 52.480 28.725 ;
        RECT 49.620 28.355 52.485 28.720 ;
        RECT 57.600 28.700 57.980 28.725 ;
        RECT 57.585 28.380 59.730 28.700 ;
        RECT 52.100 28.345 52.480 28.355 ;
        RECT 57.600 28.345 57.980 28.380 ;
        RECT 60.645 28.345 61.980 28.725 ;
        RECT 65.600 28.705 65.980 28.725 ;
        RECT 63.135 28.385 66.045 28.705 ;
        RECT 82.800 28.680 83.180 28.715 ;
        RECT 65.600 28.345 65.980 28.385 ;
        RECT 82.535 28.370 85.545 28.680 ;
        RECT 82.800 28.335 83.180 28.370 ;
        RECT 86.800 28.335 87.890 28.715 ;
        RECT 90.800 28.710 91.180 28.715 ;
        RECT 88.320 28.345 91.185 28.710 ;
        RECT 96.300 28.690 96.680 28.715 ;
        RECT 96.285 28.370 98.430 28.690 ;
        RECT 90.800 28.335 91.180 28.345 ;
        RECT 96.300 28.335 96.680 28.370 ;
        RECT 99.345 28.335 100.680 28.715 ;
        RECT 104.300 28.695 104.680 28.715 ;
        RECT 101.835 28.375 104.745 28.695 ;
        RECT 104.300 28.335 104.680 28.375 ;
        RECT 108.930 28.195 109.310 28.575 ;
        RECT 111.335 28.210 113.115 28.500 ;
        RECT 114.590 28.300 115.780 28.585 ;
        RECT 118.710 28.180 120.020 28.500 ;
        RECT 124.390 28.195 124.770 28.575 ;
        RECT 130.050 28.300 131.240 28.585 ;
        RECT 11.810 27.605 12.190 27.985 ;
        RECT 18.265 27.635 18.645 28.015 ;
        RECT 27.270 27.605 27.650 27.985 ;
        RECT 31.015 27.645 31.395 28.025 ;
        RECT 33.725 27.635 34.105 28.015 ;
        RECT 35.135 27.480 38.315 27.800 ;
        RECT 110.065 27.595 110.445 27.975 ;
        RECT 113.810 27.635 114.190 28.015 ;
        RECT 116.520 27.625 116.900 28.005 ;
        RECT 117.930 27.470 121.110 27.790 ;
        RECT 129.270 27.635 129.650 28.015 ;
        RECT 133.390 27.470 136.570 27.790 ;
        RECT 44.640 27.035 45.925 27.415 ;
        RECT 63.955 27.035 65.440 27.415 ;
        RECT 81.150 27.025 82.640 27.405 ;
        RECT 104.840 27.025 105.915 27.405 ;
        RECT 44.100 26.345 45.190 26.725 ;
        RECT 48.585 26.350 61.435 26.685 ;
        RECT 65.600 26.680 65.980 26.725 ;
        RECT 64.865 26.380 66.175 26.680 ;
        RECT 65.600 26.345 65.980 26.380 ;
        RECT 82.800 26.335 83.890 26.715 ;
        RECT 87.285 26.340 100.135 26.675 ;
        RECT 104.300 26.670 104.680 26.715 ;
        RECT 103.565 26.370 104.875 26.670 ;
        RECT 123.670 26.385 127.820 26.655 ;
        RECT 104.300 26.335 104.680 26.370 ;
        RECT 73.360 25.835 106.310 25.840 ;
        RECT 40.955 25.485 106.310 25.835 ;
        RECT 73.360 25.475 106.310 25.485 ;
        RECT 108.105 25.465 112.365 25.820 ;
        RECT 75.825 13.630 93.150 13.930 ;
        RECT 75.585 12.885 93.150 13.185 ;
        RECT 80.865 10.975 84.995 11.275 ;
        RECT 87.370 10.925 91.870 11.235 ;
        RECT 82.095 9.210 85.015 9.510 ;
        RECT 88.560 9.195 91.930 9.495 ;
      LAYER Metal2 ;
        RECT 11.950 323.970 12.250 330.900 ;
        RECT 13.260 324.570 13.560 330.920 ;
        RECT 14.575 324.600 14.870 331.425 ;
        RECT 18.415 323.970 18.715 330.910 ;
        RECT 20.625 324.545 20.930 330.905 ;
        RECT 21.475 324.545 21.775 331.365 ;
        RECT 23.285 327.990 23.665 328.370 ;
        RECT 23.500 323.280 23.880 326.300 ;
        RECT 27.410 323.970 27.710 330.900 ;
        RECT 28.720 324.570 29.020 330.920 ;
        RECT 30.035 324.600 30.330 331.425 ;
        RECT 33.875 323.970 34.175 330.910 ;
        RECT 36.085 324.545 36.405 330.905 ;
        RECT 36.935 324.545 37.235 331.365 ;
        RECT 38.710 325.945 39.090 326.325 ;
        RECT 39.415 321.830 39.775 328.390 ;
        RECT 40.555 326.580 40.880 328.445 ;
        RECT 41.220 323.235 41.680 327.920 ;
        RECT 42.005 325.780 42.455 334.600 ;
        RECT 44.190 327.605 44.620 330.595 ;
        RECT 41.935 321.890 42.315 322.270 ;
        RECT 44.825 321.910 45.205 323.285 ;
        RECT 45.595 322.730 45.910 333.780 ;
        RECT 46.610 332.475 46.900 334.535 ;
        RECT 46.530 324.620 46.855 326.990 ;
        RECT 48.180 326.665 48.580 330.630 ;
        RECT 48.900 322.560 49.225 325.325 ;
        RECT 49.885 324.595 50.290 327.925 ;
        RECT 54.535 321.620 54.905 330.720 ;
        RECT 55.480 322.685 55.770 334.520 ;
        RECT 63.385 332.415 63.695 334.930 ;
        RECT 59.295 324.650 59.735 327.925 ;
        RECT 61.675 326.665 62.200 330.605 ;
        RECT 60.835 322.560 61.160 325.325 ;
        RECT 63.350 324.655 63.765 327.045 ;
        RECT 64.380 323.215 64.695 333.900 ;
        RECT 65.710 327.605 66.195 330.615 ;
        RECT 65.080 321.825 65.415 323.175 ;
        RECT 4.795 306.000 5.150 319.790 ;
        RECT 68.140 319.160 68.590 329.425 ;
        RECT 6.420 306.855 6.780 318.190 ;
        RECT 69.305 317.620 69.790 326.505 ;
        RECT 75.610 317.245 76.015 328.775 ;
        RECT 77.685 319.145 78.075 330.245 ;
        RECT 81.455 322.695 81.810 333.780 ;
        RECT 85.200 332.420 85.490 334.480 ;
        RECT 91.980 331.270 92.290 331.300 ;
        RECT 82.780 327.550 83.250 330.540 ;
        RECT 85.130 324.565 85.445 326.935 ;
        RECT 86.750 326.610 87.170 330.575 ;
        RECT 83.415 321.855 83.795 323.230 ;
        RECT 87.490 322.505 87.815 325.270 ;
        RECT 88.475 324.540 88.880 327.870 ;
        RECT 91.980 325.170 92.295 331.270 ;
        RECT 93.125 321.565 93.495 330.665 ;
        RECT 94.070 322.630 94.360 334.465 ;
        RECT 101.975 332.360 102.285 334.875 ;
        RECT 106.225 334.060 106.605 334.440 ;
        RECT 108.355 334.060 108.735 334.440 ;
        RECT 94.965 325.125 95.295 331.320 ;
        RECT 97.870 324.595 98.325 327.870 ;
        RECT 100.230 326.610 100.775 330.550 ;
        RECT 104.285 327.550 104.720 330.560 ;
        RECT 99.425 322.505 99.750 325.270 ;
        RECT 101.940 324.600 102.355 326.990 ;
        RECT 105.480 323.175 105.810 333.870 ;
        RECT 106.915 327.510 107.300 333.295 ;
        RECT 103.670 321.770 104.005 323.120 ;
        RECT 107.275 322.755 107.700 327.030 ;
        RECT 108.975 324.520 109.275 331.560 ;
        RECT 105.935 321.845 106.315 322.225 ;
        RECT 108.130 321.830 108.510 322.210 ;
        RECT 112.000 321.770 112.290 331.550 ;
        RECT 113.850 324.005 114.150 330.815 ;
        RECT 114.640 324.600 114.950 334.640 ;
        RECT 123.830 332.885 124.210 333.265 ;
        RECT 115.435 324.530 115.735 331.360 ;
        RECT 118.010 323.790 118.290 326.825 ;
        RECT 120.760 323.745 121.060 330.900 ;
        RECT 124.435 324.520 124.735 331.560 ;
        RECT 123.730 322.710 124.110 323.090 ;
        RECT 127.460 322.305 127.750 331.550 ;
        RECT 129.310 324.005 129.610 330.815 ;
        RECT 130.100 324.600 130.410 333.335 ;
        RECT 130.895 324.530 131.195 331.360 ;
        RECT 133.470 323.790 133.750 326.825 ;
        RECT 136.220 323.745 136.520 330.900 ;
        RECT 11.905 304.280 12.205 311.210 ;
        RECT 13.215 304.880 13.515 311.230 ;
        RECT 14.530 304.910 14.825 311.735 ;
        RECT 18.370 304.280 18.670 311.220 ;
        RECT 20.580 304.855 20.885 311.215 ;
        RECT 21.430 304.855 21.730 311.675 ;
        RECT 23.240 308.300 23.620 308.680 ;
        RECT 25.025 306.880 25.345 309.010 ;
        RECT 23.455 303.590 23.835 306.610 ;
        RECT 25.635 306.040 25.915 308.445 ;
        RECT 26.245 304.885 26.545 311.925 ;
        RECT 27.365 304.280 27.665 311.210 ;
        RECT 28.675 304.880 28.975 311.230 ;
        RECT 29.270 306.755 29.595 311.915 ;
        RECT 29.990 304.910 30.285 311.735 ;
        RECT 31.120 304.370 31.420 311.180 ;
        RECT 31.910 304.965 32.220 311.155 ;
        RECT 32.705 304.895 33.005 311.725 ;
        RECT 33.830 304.280 34.130 311.220 ;
        RECT 35.280 304.155 35.560 307.190 ;
        RECT 36.040 304.855 36.360 311.215 ;
        RECT 36.890 304.855 37.190 311.675 ;
        RECT 38.030 304.110 38.330 311.265 ;
        RECT 38.665 306.255 39.045 306.635 ;
        RECT 39.370 302.140 39.730 308.700 ;
        RECT 40.510 306.890 40.835 308.755 ;
        RECT 41.175 303.545 41.635 308.230 ;
        RECT 41.960 306.090 42.410 314.910 ;
        RECT 44.145 307.915 44.575 310.905 ;
        RECT 41.890 302.200 42.270 302.580 ;
        RECT 44.780 302.220 45.160 303.595 ;
        RECT 45.550 303.040 45.865 314.090 ;
        RECT 46.565 312.785 46.855 314.845 ;
        RECT 46.485 304.930 46.810 307.300 ;
        RECT 48.135 306.975 48.535 310.940 ;
        RECT 48.855 302.870 49.180 305.635 ;
        RECT 49.840 304.905 50.245 308.235 ;
        RECT 54.490 301.930 54.860 311.030 ;
        RECT 55.435 302.995 55.725 314.830 ;
        RECT 63.340 312.725 63.650 315.240 ;
        RECT 59.250 304.960 59.690 308.235 ;
        RECT 61.630 306.975 62.155 310.915 ;
        RECT 60.790 302.870 61.115 305.635 ;
        RECT 63.305 304.965 63.720 307.355 ;
        RECT 64.335 303.525 64.650 314.210 ;
        RECT 65.665 307.915 66.150 310.925 ;
        RECT 65.035 302.135 65.370 303.485 ;
        RECT 4.795 286.235 5.150 300.290 ;
        RECT 68.140 299.660 68.590 309.775 ;
        RECT 6.420 287.040 6.780 298.690 ;
        RECT 69.305 298.120 69.790 306.875 ;
        RECT 75.910 297.495 76.315 309.025 ;
        RECT 77.985 299.395 78.375 310.495 ;
        RECT 81.255 302.970 81.610 314.055 ;
        RECT 85.000 312.695 85.290 314.755 ;
        RECT 91.780 311.545 92.090 311.575 ;
        RECT 82.580 307.825 83.050 310.815 ;
        RECT 84.930 304.840 85.245 307.210 ;
        RECT 86.550 306.885 86.970 310.850 ;
        RECT 83.215 302.130 83.595 303.505 ;
        RECT 87.290 302.780 87.615 305.545 ;
        RECT 88.275 304.815 88.680 308.145 ;
        RECT 91.780 305.445 92.095 311.545 ;
        RECT 92.925 301.840 93.295 310.940 ;
        RECT 93.870 302.905 94.160 314.740 ;
        RECT 101.775 312.635 102.085 315.150 ;
        RECT 106.025 314.335 106.405 314.715 ;
        RECT 108.155 314.335 108.535 314.715 ;
        RECT 94.765 305.400 95.095 311.595 ;
        RECT 97.670 304.870 98.125 308.145 ;
        RECT 100.030 306.885 100.575 310.825 ;
        RECT 104.085 307.825 104.520 310.835 ;
        RECT 99.225 302.780 99.550 305.545 ;
        RECT 101.740 304.875 102.155 307.265 ;
        RECT 105.280 303.450 105.610 314.145 ;
        RECT 106.715 307.785 107.100 313.570 ;
        RECT 103.470 302.045 103.805 303.395 ;
        RECT 107.075 303.030 107.500 307.305 ;
        RECT 108.775 304.795 109.075 311.835 ;
        RECT 109.895 304.190 110.195 311.120 ;
        RECT 111.205 304.790 111.505 311.140 ;
        RECT 105.735 302.120 106.115 302.500 ;
        RECT 107.930 302.105 108.310 302.485 ;
        RECT 111.800 302.045 112.090 311.825 ;
        RECT 112.520 304.820 112.815 311.645 ;
        RECT 113.650 304.280 113.950 311.090 ;
        RECT 114.440 304.875 114.750 314.915 ;
        RECT 123.630 313.160 124.010 313.540 ;
        RECT 115.235 304.805 115.535 311.635 ;
        RECT 116.360 304.190 116.660 311.130 ;
        RECT 117.810 304.065 118.090 307.100 ;
        RECT 118.570 304.765 118.850 311.125 ;
        RECT 119.420 304.765 119.720 311.585 ;
        RECT 120.560 304.020 120.860 311.175 ;
        RECT 121.205 308.210 121.585 308.590 ;
        RECT 121.205 306.155 121.585 306.535 ;
        RECT 123.055 306.035 123.370 310.360 ;
        RECT 123.665 308.110 123.945 309.640 ;
        RECT 124.235 304.795 124.535 311.835 ;
        RECT 126.010 305.550 126.310 309.610 ;
        RECT 123.530 302.985 123.910 303.365 ;
        RECT 127.260 302.580 127.550 311.825 ;
        RECT 129.110 304.280 129.410 311.090 ;
        RECT 129.900 304.875 130.210 313.610 ;
        RECT 130.695 304.805 130.995 311.635 ;
        RECT 132.500 305.535 132.780 309.625 ;
        RECT 133.270 304.065 133.550 307.100 ;
        RECT 136.020 304.020 136.320 311.175 ;
        RECT 138.060 309.915 138.435 318.115 ;
        RECT 139.805 309.110 140.105 320.105 ;
        RECT 12.095 284.570 12.395 291.500 ;
        RECT 13.405 285.170 13.705 291.520 ;
        RECT 14.720 285.200 15.015 292.025 ;
        RECT 18.560 284.570 18.860 291.510 ;
        RECT 20.770 285.145 21.075 291.505 ;
        RECT 21.620 285.145 21.920 291.965 ;
        RECT 23.430 288.590 23.810 288.970 ;
        RECT 25.215 287.170 25.535 289.300 ;
        RECT 23.645 283.880 24.025 286.900 ;
        RECT 25.825 286.330 26.105 288.735 ;
        RECT 26.435 285.175 26.735 292.215 ;
        RECT 27.555 284.570 27.855 291.500 ;
        RECT 28.865 285.170 29.165 291.520 ;
        RECT 29.460 287.045 29.785 292.205 ;
        RECT 30.180 285.200 30.475 292.025 ;
        RECT 31.310 284.660 31.610 291.470 ;
        RECT 32.100 285.255 32.410 291.445 ;
        RECT 32.895 285.185 33.195 292.015 ;
        RECT 34.020 284.570 34.320 291.510 ;
        RECT 35.470 284.445 35.750 287.480 ;
        RECT 36.230 285.145 36.550 291.505 ;
        RECT 37.080 285.145 37.380 291.965 ;
        RECT 38.220 284.400 38.520 291.555 ;
        RECT 38.855 286.545 39.235 286.925 ;
        RECT 39.560 282.430 39.920 288.990 ;
        RECT 40.700 287.180 41.025 289.045 ;
        RECT 41.365 283.835 41.825 288.520 ;
        RECT 42.150 286.380 42.600 295.200 ;
        RECT 44.335 288.205 44.765 291.195 ;
        RECT 42.080 282.490 42.460 282.870 ;
        RECT 44.970 282.510 45.350 283.885 ;
        RECT 45.740 283.330 46.055 294.380 ;
        RECT 46.755 293.075 47.045 295.135 ;
        RECT 46.675 285.220 47.000 287.590 ;
        RECT 48.325 287.265 48.725 291.230 ;
        RECT 49.045 283.160 49.370 285.925 ;
        RECT 50.030 285.195 50.435 288.525 ;
        RECT 54.680 282.220 55.050 291.320 ;
        RECT 55.625 283.285 55.915 295.120 ;
        RECT 63.530 293.015 63.840 295.530 ;
        RECT 59.440 285.250 59.880 288.525 ;
        RECT 61.820 287.265 62.345 291.205 ;
        RECT 60.980 283.160 61.305 285.925 ;
        RECT 63.495 285.255 63.910 287.645 ;
        RECT 64.525 283.815 64.840 294.500 ;
        RECT 65.855 288.205 66.340 291.215 ;
        RECT 65.225 282.425 65.560 283.775 ;
        RECT 5.005 266.460 5.360 280.250 ;
        RECT 68.350 279.620 68.800 290.120 ;
        RECT 6.630 267.315 6.990 278.650 ;
        RECT 69.515 278.080 70.000 287.320 ;
        RECT 75.930 277.835 76.335 289.365 ;
        RECT 78.005 279.735 78.395 290.835 ;
        RECT 81.410 283.325 81.765 294.410 ;
        RECT 85.155 293.050 85.445 295.110 ;
        RECT 91.935 291.900 92.245 291.930 ;
        RECT 82.735 288.180 83.205 291.170 ;
        RECT 85.085 285.195 85.400 287.565 ;
        RECT 86.705 287.240 87.125 291.205 ;
        RECT 83.370 282.485 83.750 283.860 ;
        RECT 87.445 283.135 87.770 285.900 ;
        RECT 88.430 285.170 88.835 288.500 ;
        RECT 91.935 285.800 92.250 291.900 ;
        RECT 93.080 282.195 93.450 291.295 ;
        RECT 94.025 283.260 94.315 295.095 ;
        RECT 101.930 292.990 102.240 295.505 ;
        RECT 106.180 294.690 106.560 295.070 ;
        RECT 108.310 294.690 108.690 295.070 ;
        RECT 94.920 285.755 95.250 291.950 ;
        RECT 97.825 285.225 98.280 288.500 ;
        RECT 100.185 287.240 100.730 291.180 ;
        RECT 104.240 288.180 104.675 291.190 ;
        RECT 99.380 283.135 99.705 285.900 ;
        RECT 101.895 285.230 102.310 287.620 ;
        RECT 105.435 283.805 105.765 294.500 ;
        RECT 106.870 288.140 107.255 293.925 ;
        RECT 103.625 282.400 103.960 283.750 ;
        RECT 107.230 283.385 107.655 287.660 ;
        RECT 108.930 285.150 109.230 292.190 ;
        RECT 110.050 284.545 110.350 291.475 ;
        RECT 111.360 285.145 111.660 291.495 ;
        RECT 105.890 282.475 106.270 282.855 ;
        RECT 108.085 282.460 108.465 282.840 ;
        RECT 111.955 282.400 112.245 292.180 ;
        RECT 112.675 285.175 112.970 292.000 ;
        RECT 113.805 284.635 114.105 291.445 ;
        RECT 114.595 285.230 114.905 295.270 ;
        RECT 123.785 293.515 124.165 293.895 ;
        RECT 115.390 285.160 115.690 291.990 ;
        RECT 116.515 284.545 116.815 291.485 ;
        RECT 117.965 284.420 118.245 287.455 ;
        RECT 118.725 285.120 119.005 291.480 ;
        RECT 119.575 285.120 119.875 291.940 ;
        RECT 120.715 284.375 121.015 291.530 ;
        RECT 121.360 288.565 121.740 288.945 ;
        RECT 121.360 286.510 121.740 286.890 ;
        RECT 123.210 286.390 123.525 290.715 ;
        RECT 123.820 288.465 124.100 289.995 ;
        RECT 124.390 285.150 124.690 292.190 ;
        RECT 126.165 285.905 126.465 289.965 ;
        RECT 123.685 283.340 124.065 283.720 ;
        RECT 127.415 282.935 127.705 292.180 ;
        RECT 129.265 284.635 129.565 291.445 ;
        RECT 130.055 285.230 130.365 293.965 ;
        RECT 130.850 285.160 131.150 291.990 ;
        RECT 132.655 285.890 132.935 289.980 ;
        RECT 133.425 284.420 133.705 287.455 ;
        RECT 136.175 284.375 136.475 291.530 ;
        RECT 138.360 290.165 138.735 298.365 ;
        RECT 140.105 289.360 140.405 300.355 ;
        RECT 11.900 264.730 12.200 271.660 ;
        RECT 13.210 265.330 13.510 271.680 ;
        RECT 14.525 265.360 14.820 272.185 ;
        RECT 18.365 264.730 18.665 271.670 ;
        RECT 20.575 265.305 20.880 271.665 ;
        RECT 21.425 265.305 21.725 272.125 ;
        RECT 23.235 268.750 23.615 269.130 ;
        RECT 25.020 267.330 25.340 269.460 ;
        RECT 23.450 264.040 23.830 267.060 ;
        RECT 25.630 266.490 25.910 268.895 ;
        RECT 26.240 265.335 26.540 272.375 ;
        RECT 27.360 264.730 27.660 271.660 ;
        RECT 28.670 265.330 28.970 271.680 ;
        RECT 29.265 267.205 29.590 272.365 ;
        RECT 29.985 265.360 30.280 272.185 ;
        RECT 31.115 264.820 31.415 271.630 ;
        RECT 31.905 265.415 32.215 271.605 ;
        RECT 32.700 265.345 33.000 272.175 ;
        RECT 33.825 264.730 34.125 271.670 ;
        RECT 35.275 264.605 35.555 267.640 ;
        RECT 36.035 265.305 36.355 271.665 ;
        RECT 36.885 265.305 37.185 272.125 ;
        RECT 38.025 264.560 38.325 271.715 ;
        RECT 38.660 266.705 39.040 267.085 ;
        RECT 39.365 262.590 39.725 269.150 ;
        RECT 40.505 267.340 40.830 269.205 ;
        RECT 41.170 263.995 41.630 268.680 ;
        RECT 41.955 266.540 42.405 275.360 ;
        RECT 44.140 268.365 44.570 271.355 ;
        RECT 41.885 262.650 42.265 263.030 ;
        RECT 44.775 262.670 45.155 264.045 ;
        RECT 45.545 263.490 45.860 274.540 ;
        RECT 46.560 273.235 46.850 275.295 ;
        RECT 46.480 265.380 46.805 267.750 ;
        RECT 48.130 267.425 48.530 271.390 ;
        RECT 48.850 263.320 49.175 266.085 ;
        RECT 49.835 265.355 50.240 268.685 ;
        RECT 54.485 262.380 54.855 271.480 ;
        RECT 55.430 263.445 55.720 275.280 ;
        RECT 63.335 273.175 63.645 275.690 ;
        RECT 59.245 265.410 59.685 268.685 ;
        RECT 61.625 267.425 62.150 271.365 ;
        RECT 60.785 263.320 61.110 266.085 ;
        RECT 63.300 265.415 63.715 267.805 ;
        RECT 64.330 263.975 64.645 274.660 ;
        RECT 65.660 268.365 66.145 271.375 ;
        RECT 65.030 262.585 65.365 263.935 ;
        RECT 4.960 246.670 5.315 260.460 ;
        RECT 68.305 259.830 68.755 270.320 ;
        RECT 6.585 247.575 6.945 258.860 ;
        RECT 69.470 258.290 69.955 267.450 ;
        RECT 75.930 258.100 76.335 269.630 ;
        RECT 78.005 260.000 78.395 271.100 ;
        RECT 81.410 263.530 81.765 274.615 ;
        RECT 85.155 273.255 85.445 275.315 ;
        RECT 91.935 272.105 92.245 272.135 ;
        RECT 82.735 268.385 83.205 271.375 ;
        RECT 85.085 265.400 85.400 267.770 ;
        RECT 86.705 267.445 87.125 271.410 ;
        RECT 83.370 262.690 83.750 264.065 ;
        RECT 87.445 263.340 87.770 266.105 ;
        RECT 88.430 265.375 88.835 268.705 ;
        RECT 91.935 266.005 92.250 272.105 ;
        RECT 93.080 262.400 93.450 271.500 ;
        RECT 94.025 263.465 94.315 275.300 ;
        RECT 101.930 273.195 102.240 275.710 ;
        RECT 106.180 274.895 106.560 275.275 ;
        RECT 108.310 274.895 108.690 275.275 ;
        RECT 94.920 265.960 95.250 272.155 ;
        RECT 97.825 265.430 98.280 268.705 ;
        RECT 100.185 267.445 100.730 271.385 ;
        RECT 104.240 268.385 104.675 271.395 ;
        RECT 99.380 263.340 99.705 266.105 ;
        RECT 101.895 265.435 102.310 267.825 ;
        RECT 105.435 264.010 105.765 274.705 ;
        RECT 106.870 268.345 107.255 274.130 ;
        RECT 103.625 262.605 103.960 263.955 ;
        RECT 107.230 263.590 107.655 267.865 ;
        RECT 108.930 265.355 109.230 272.395 ;
        RECT 110.050 264.750 110.350 271.680 ;
        RECT 111.360 265.350 111.660 271.700 ;
        RECT 105.890 262.680 106.270 263.060 ;
        RECT 108.085 262.665 108.465 263.045 ;
        RECT 111.955 262.605 112.245 272.385 ;
        RECT 112.675 265.380 112.970 272.205 ;
        RECT 113.805 264.840 114.105 271.650 ;
        RECT 114.595 265.435 114.905 275.475 ;
        RECT 123.785 273.720 124.165 274.100 ;
        RECT 115.390 265.365 115.690 272.195 ;
        RECT 116.515 264.750 116.815 271.690 ;
        RECT 117.965 264.625 118.245 267.660 ;
        RECT 118.725 265.325 119.005 271.685 ;
        RECT 119.575 265.325 119.875 272.145 ;
        RECT 120.715 264.580 121.015 271.735 ;
        RECT 121.360 268.770 121.740 269.150 ;
        RECT 121.360 266.715 121.740 267.095 ;
        RECT 123.210 266.595 123.525 270.920 ;
        RECT 123.820 268.670 124.100 270.200 ;
        RECT 124.390 265.355 124.690 272.395 ;
        RECT 126.165 266.110 126.465 270.170 ;
        RECT 123.685 263.545 124.065 263.925 ;
        RECT 127.415 263.140 127.705 272.385 ;
        RECT 129.265 264.840 129.565 271.650 ;
        RECT 130.055 265.435 130.365 274.170 ;
        RECT 130.850 265.365 131.150 272.195 ;
        RECT 132.655 266.095 132.935 270.185 ;
        RECT 133.425 264.625 133.705 267.660 ;
        RECT 136.175 264.580 136.475 271.735 ;
        RECT 138.380 270.505 138.755 278.705 ;
        RECT 140.125 269.700 140.425 280.695 ;
        RECT 11.770 245.020 12.070 251.950 ;
        RECT 13.080 245.620 13.380 251.970 ;
        RECT 14.395 245.650 14.690 252.475 ;
        RECT 18.235 245.020 18.535 251.960 ;
        RECT 20.445 245.595 20.750 251.955 ;
        RECT 21.295 245.595 21.595 252.415 ;
        RECT 23.105 249.040 23.485 249.420 ;
        RECT 24.890 247.620 25.210 249.750 ;
        RECT 23.320 244.330 23.700 247.350 ;
        RECT 25.500 246.780 25.780 249.185 ;
        RECT 26.110 245.625 26.410 252.665 ;
        RECT 27.230 245.020 27.530 251.950 ;
        RECT 28.540 245.620 28.840 251.970 ;
        RECT 29.135 247.495 29.460 252.655 ;
        RECT 29.855 245.650 30.150 252.475 ;
        RECT 30.985 245.110 31.285 251.920 ;
        RECT 31.775 245.705 32.085 251.895 ;
        RECT 32.570 245.635 32.870 252.465 ;
        RECT 33.695 245.020 33.995 251.960 ;
        RECT 35.145 244.895 35.425 247.930 ;
        RECT 35.905 245.595 36.225 251.955 ;
        RECT 36.755 245.595 37.055 252.415 ;
        RECT 37.895 244.850 38.195 252.005 ;
        RECT 38.530 246.995 38.910 247.375 ;
        RECT 39.235 242.880 39.595 249.440 ;
        RECT 40.375 247.630 40.700 249.495 ;
        RECT 41.040 244.285 41.500 248.970 ;
        RECT 41.825 246.830 42.275 255.650 ;
        RECT 44.010 248.655 44.440 251.645 ;
        RECT 41.755 242.940 42.135 243.320 ;
        RECT 44.645 242.960 45.025 244.335 ;
        RECT 45.415 243.780 45.730 254.830 ;
        RECT 46.430 253.525 46.720 255.585 ;
        RECT 46.350 245.670 46.675 248.040 ;
        RECT 48.000 247.715 48.400 251.680 ;
        RECT 48.720 243.610 49.045 246.375 ;
        RECT 49.705 245.645 50.110 248.975 ;
        RECT 54.355 242.670 54.725 251.770 ;
        RECT 55.300 243.735 55.590 255.570 ;
        RECT 63.205 253.465 63.515 255.980 ;
        RECT 59.115 245.700 59.555 248.975 ;
        RECT 61.495 247.715 62.020 251.655 ;
        RECT 60.655 243.610 60.980 246.375 ;
        RECT 63.170 245.705 63.585 248.095 ;
        RECT 64.200 244.265 64.515 254.950 ;
        RECT 65.530 248.655 66.015 251.665 ;
        RECT 64.900 242.875 65.235 244.225 ;
        RECT 4.655 226.910 5.010 240.830 ;
        RECT 68.000 240.200 68.450 250.465 ;
        RECT 6.280 227.815 6.640 239.230 ;
        RECT 69.165 238.660 69.650 247.545 ;
        RECT 75.830 238.395 76.235 249.925 ;
        RECT 77.905 240.295 78.295 251.395 ;
        RECT 81.330 243.775 81.685 254.860 ;
        RECT 85.075 253.500 85.365 255.560 ;
        RECT 91.855 252.350 92.165 252.380 ;
        RECT 82.655 248.630 83.125 251.620 ;
        RECT 85.005 245.645 85.320 248.015 ;
        RECT 86.625 247.690 87.045 251.655 ;
        RECT 83.290 242.935 83.670 244.310 ;
        RECT 87.365 243.585 87.690 246.350 ;
        RECT 88.350 245.620 88.755 248.950 ;
        RECT 91.855 246.250 92.170 252.350 ;
        RECT 93.000 242.645 93.370 251.745 ;
        RECT 93.945 243.710 94.235 255.545 ;
        RECT 101.850 253.440 102.160 255.955 ;
        RECT 106.100 255.140 106.480 255.520 ;
        RECT 108.230 255.140 108.610 255.520 ;
        RECT 94.840 246.205 95.170 252.400 ;
        RECT 97.745 245.675 98.200 248.950 ;
        RECT 100.105 247.690 100.650 251.630 ;
        RECT 104.160 248.630 104.595 251.640 ;
        RECT 99.300 243.585 99.625 246.350 ;
        RECT 101.815 245.680 102.230 248.070 ;
        RECT 105.355 244.255 105.685 254.950 ;
        RECT 106.790 248.590 107.175 254.375 ;
        RECT 103.545 242.850 103.880 244.200 ;
        RECT 107.150 243.835 107.575 248.110 ;
        RECT 108.850 245.600 109.150 252.640 ;
        RECT 109.970 244.995 110.270 251.925 ;
        RECT 111.280 245.595 111.580 251.945 ;
        RECT 105.810 242.925 106.190 243.305 ;
        RECT 108.005 242.910 108.385 243.290 ;
        RECT 111.875 242.850 112.165 252.630 ;
        RECT 112.595 245.625 112.890 252.450 ;
        RECT 113.725 245.085 114.025 251.895 ;
        RECT 114.515 245.680 114.825 255.720 ;
        RECT 123.705 253.965 124.085 254.345 ;
        RECT 115.310 245.610 115.610 252.440 ;
        RECT 116.435 244.995 116.735 251.935 ;
        RECT 117.885 244.870 118.165 247.905 ;
        RECT 118.645 245.570 118.925 251.930 ;
        RECT 119.495 245.570 119.795 252.390 ;
        RECT 120.635 244.825 120.935 251.980 ;
        RECT 121.280 249.015 121.660 249.395 ;
        RECT 121.280 246.960 121.660 247.340 ;
        RECT 123.130 246.840 123.445 251.165 ;
        RECT 123.740 248.915 124.020 250.445 ;
        RECT 124.310 245.600 124.610 252.640 ;
        RECT 126.085 246.355 126.385 250.415 ;
        RECT 123.605 243.790 123.985 244.170 ;
        RECT 127.335 243.385 127.625 252.630 ;
        RECT 129.185 245.085 129.485 251.895 ;
        RECT 129.975 245.680 130.285 254.415 ;
        RECT 130.770 245.610 131.070 252.440 ;
        RECT 132.575 246.340 132.855 250.430 ;
        RECT 133.345 244.870 133.625 247.905 ;
        RECT 136.095 244.825 136.395 251.980 ;
        RECT 138.380 250.685 138.755 258.970 ;
        RECT 140.125 249.965 140.425 260.960 ;
        RECT 11.900 225.260 12.200 232.190 ;
        RECT 13.210 225.860 13.510 232.210 ;
        RECT 14.525 225.890 14.820 232.715 ;
        RECT 18.365 225.260 18.665 232.200 ;
        RECT 20.575 225.835 20.880 232.195 ;
        RECT 21.425 225.835 21.725 232.655 ;
        RECT 23.235 229.280 23.615 229.660 ;
        RECT 25.020 227.860 25.340 229.990 ;
        RECT 23.450 224.570 23.830 227.590 ;
        RECT 25.630 227.020 25.910 229.425 ;
        RECT 26.240 225.865 26.540 232.905 ;
        RECT 27.360 225.260 27.660 232.190 ;
        RECT 28.670 225.860 28.970 232.210 ;
        RECT 29.265 227.735 29.590 232.895 ;
        RECT 29.985 225.890 30.280 232.715 ;
        RECT 31.115 225.350 31.415 232.160 ;
        RECT 31.905 225.945 32.215 232.135 ;
        RECT 32.700 225.875 33.000 232.705 ;
        RECT 33.825 225.260 34.125 232.200 ;
        RECT 35.275 225.135 35.555 228.170 ;
        RECT 36.035 225.835 36.355 232.195 ;
        RECT 36.885 225.835 37.185 232.655 ;
        RECT 38.025 225.090 38.325 232.245 ;
        RECT 38.660 227.235 39.040 227.615 ;
        RECT 39.365 223.120 39.725 229.680 ;
        RECT 40.505 227.870 40.830 229.735 ;
        RECT 41.170 224.525 41.630 229.210 ;
        RECT 41.955 227.070 42.405 235.890 ;
        RECT 44.140 228.895 44.570 231.885 ;
        RECT 41.885 223.180 42.265 223.560 ;
        RECT 44.775 223.200 45.155 224.575 ;
        RECT 45.545 224.020 45.860 235.070 ;
        RECT 46.560 233.765 46.850 235.825 ;
        RECT 46.480 225.910 46.805 228.280 ;
        RECT 48.130 227.955 48.530 231.920 ;
        RECT 48.850 223.850 49.175 226.615 ;
        RECT 49.835 225.885 50.240 229.215 ;
        RECT 54.485 222.910 54.855 232.010 ;
        RECT 55.430 223.975 55.720 235.810 ;
        RECT 63.335 233.705 63.645 236.220 ;
        RECT 59.245 225.940 59.685 229.215 ;
        RECT 61.625 227.955 62.150 231.895 ;
        RECT 60.785 223.850 61.110 226.615 ;
        RECT 63.300 225.945 63.715 228.335 ;
        RECT 64.330 224.505 64.645 235.190 ;
        RECT 65.660 228.895 66.145 231.905 ;
        RECT 65.030 223.115 65.365 224.465 ;
        RECT 4.750 207.145 5.105 221.055 ;
        RECT 68.095 220.425 68.545 230.690 ;
        RECT 6.375 208.065 6.735 219.455 ;
        RECT 69.260 218.885 69.745 227.770 ;
        RECT 76.090 218.240 76.495 230.120 ;
        RECT 78.165 220.140 78.555 231.720 ;
        RECT 81.435 224.060 81.790 235.145 ;
        RECT 85.180 233.785 85.470 235.845 ;
        RECT 91.960 232.635 92.270 232.665 ;
        RECT 82.760 228.915 83.230 231.905 ;
        RECT 85.110 225.930 85.425 228.300 ;
        RECT 86.730 227.975 87.150 231.940 ;
        RECT 83.395 223.220 83.775 224.595 ;
        RECT 87.470 223.870 87.795 226.635 ;
        RECT 88.455 225.905 88.860 229.235 ;
        RECT 91.960 226.535 92.275 232.635 ;
        RECT 93.105 222.930 93.475 232.030 ;
        RECT 94.050 223.995 94.340 235.830 ;
        RECT 101.955 233.725 102.265 236.240 ;
        RECT 106.205 235.425 106.585 235.805 ;
        RECT 108.335 235.425 108.715 235.805 ;
        RECT 94.945 226.490 95.275 232.685 ;
        RECT 97.850 225.960 98.305 229.235 ;
        RECT 100.210 227.975 100.755 231.915 ;
        RECT 104.265 228.915 104.700 231.925 ;
        RECT 99.405 223.870 99.730 226.635 ;
        RECT 101.920 225.965 102.335 228.355 ;
        RECT 105.460 224.540 105.790 235.235 ;
        RECT 106.895 228.875 107.280 234.660 ;
        RECT 103.650 223.135 103.985 224.485 ;
        RECT 107.255 224.120 107.680 228.395 ;
        RECT 108.955 225.885 109.255 232.925 ;
        RECT 110.075 225.280 110.375 232.210 ;
        RECT 111.385 225.880 111.685 232.230 ;
        RECT 105.915 223.210 106.295 223.590 ;
        RECT 108.110 223.195 108.490 223.575 ;
        RECT 111.980 223.135 112.270 232.915 ;
        RECT 112.700 225.910 112.995 232.735 ;
        RECT 113.830 225.370 114.130 232.180 ;
        RECT 114.620 225.965 114.930 236.005 ;
        RECT 123.810 234.250 124.190 234.630 ;
        RECT 115.415 225.895 115.715 232.725 ;
        RECT 116.540 225.280 116.840 232.220 ;
        RECT 117.990 225.155 118.270 228.190 ;
        RECT 118.750 225.855 119.030 232.215 ;
        RECT 119.600 225.855 119.900 232.675 ;
        RECT 120.740 225.110 121.040 232.265 ;
        RECT 121.385 229.300 121.765 229.680 ;
        RECT 121.385 227.245 121.765 227.625 ;
        RECT 123.235 227.125 123.550 231.450 ;
        RECT 123.845 229.200 124.125 230.730 ;
        RECT 124.415 225.885 124.715 232.925 ;
        RECT 126.190 226.640 126.490 230.700 ;
        RECT 123.710 224.075 124.090 224.455 ;
        RECT 127.440 223.670 127.730 232.915 ;
        RECT 129.290 225.370 129.590 232.180 ;
        RECT 130.080 225.965 130.390 234.700 ;
        RECT 130.875 225.895 131.175 232.725 ;
        RECT 132.680 226.625 132.960 230.715 ;
        RECT 133.450 225.155 133.730 228.190 ;
        RECT 136.200 225.110 136.500 232.265 ;
        RECT 138.280 230.985 138.655 239.265 ;
        RECT 140.025 230.145 140.325 241.255 ;
        RECT 11.850 205.450 12.150 212.380 ;
        RECT 13.160 206.050 13.460 212.400 ;
        RECT 14.475 206.080 14.770 212.905 ;
        RECT 18.315 205.450 18.615 212.390 ;
        RECT 20.525 206.025 20.830 212.385 ;
        RECT 21.375 206.025 21.675 212.845 ;
        RECT 23.185 209.470 23.565 209.850 ;
        RECT 24.970 208.050 25.290 210.180 ;
        RECT 23.400 204.760 23.780 207.780 ;
        RECT 25.580 207.210 25.860 209.615 ;
        RECT 26.190 206.055 26.490 213.095 ;
        RECT 27.310 205.450 27.610 212.380 ;
        RECT 28.620 206.050 28.920 212.400 ;
        RECT 29.215 207.925 29.540 213.085 ;
        RECT 29.935 206.080 30.230 212.905 ;
        RECT 31.065 205.540 31.365 212.350 ;
        RECT 31.855 206.135 32.165 212.325 ;
        RECT 32.650 206.065 32.950 212.895 ;
        RECT 33.775 205.450 34.075 212.390 ;
        RECT 35.225 205.325 35.505 208.360 ;
        RECT 35.985 206.025 36.305 212.385 ;
        RECT 36.835 206.025 37.135 212.845 ;
        RECT 37.975 205.280 38.275 212.435 ;
        RECT 38.610 207.425 38.990 207.805 ;
        RECT 39.315 203.310 39.675 209.870 ;
        RECT 40.455 208.060 40.780 209.925 ;
        RECT 41.120 204.715 41.580 209.400 ;
        RECT 41.905 207.260 42.355 216.080 ;
        RECT 44.090 209.085 44.520 212.075 ;
        RECT 41.835 203.370 42.215 203.750 ;
        RECT 44.725 203.390 45.105 204.765 ;
        RECT 45.495 204.210 45.810 215.260 ;
        RECT 46.510 213.955 46.800 216.015 ;
        RECT 46.430 206.100 46.755 208.470 ;
        RECT 48.080 208.145 48.480 212.110 ;
        RECT 48.800 204.040 49.125 206.805 ;
        RECT 49.785 206.075 50.190 209.405 ;
        RECT 54.435 203.100 54.805 212.200 ;
        RECT 55.380 204.165 55.670 216.000 ;
        RECT 63.285 213.895 63.595 216.410 ;
        RECT 59.195 206.130 59.635 209.405 ;
        RECT 61.575 208.145 62.100 212.085 ;
        RECT 60.735 204.040 61.060 206.805 ;
        RECT 63.250 206.135 63.665 208.525 ;
        RECT 64.280 204.695 64.595 215.380 ;
        RECT 65.610 209.085 66.095 212.095 ;
        RECT 64.980 203.305 65.315 204.655 ;
        RECT 4.750 187.305 5.105 201.245 ;
        RECT 68.095 200.615 68.545 210.880 ;
        RECT 6.375 188.095 6.735 199.645 ;
        RECT 69.260 199.075 69.745 207.960 ;
        RECT 76.200 198.350 76.605 210.395 ;
        RECT 78.275 200.250 78.665 211.675 ;
        RECT 81.435 204.090 81.790 215.175 ;
        RECT 85.180 213.815 85.470 215.875 ;
        RECT 91.960 212.665 92.270 212.695 ;
        RECT 82.760 208.945 83.230 211.935 ;
        RECT 85.110 205.960 85.425 208.330 ;
        RECT 86.730 208.005 87.150 211.970 ;
        RECT 83.395 203.250 83.775 204.625 ;
        RECT 87.470 203.900 87.795 206.665 ;
        RECT 88.455 205.935 88.860 209.265 ;
        RECT 91.960 206.565 92.275 212.665 ;
        RECT 93.105 202.960 93.475 212.060 ;
        RECT 94.050 204.025 94.340 215.860 ;
        RECT 101.955 213.755 102.265 216.270 ;
        RECT 106.205 215.455 106.585 215.835 ;
        RECT 108.335 215.455 108.715 215.835 ;
        RECT 94.945 206.520 95.275 212.715 ;
        RECT 97.850 205.990 98.305 209.265 ;
        RECT 100.210 208.005 100.755 211.945 ;
        RECT 104.265 208.945 104.700 211.955 ;
        RECT 99.405 203.900 99.730 206.665 ;
        RECT 101.920 205.995 102.335 208.385 ;
        RECT 105.460 204.570 105.790 215.265 ;
        RECT 106.895 208.905 107.280 214.690 ;
        RECT 103.650 203.165 103.985 204.515 ;
        RECT 107.255 204.150 107.680 208.425 ;
        RECT 108.955 205.915 109.255 212.955 ;
        RECT 110.075 205.310 110.375 212.240 ;
        RECT 111.385 205.910 111.685 212.260 ;
        RECT 105.915 203.240 106.295 203.620 ;
        RECT 108.110 203.225 108.490 203.605 ;
        RECT 111.980 203.165 112.270 212.945 ;
        RECT 112.700 205.940 112.995 212.765 ;
        RECT 113.830 205.400 114.130 212.210 ;
        RECT 114.620 205.995 114.930 216.035 ;
        RECT 123.810 214.280 124.190 214.660 ;
        RECT 115.415 205.925 115.715 212.755 ;
        RECT 116.540 205.310 116.840 212.250 ;
        RECT 117.990 205.185 118.270 208.220 ;
        RECT 118.750 205.885 119.030 212.245 ;
        RECT 119.600 205.885 119.900 212.705 ;
        RECT 120.740 205.140 121.040 212.295 ;
        RECT 121.385 209.330 121.765 209.710 ;
        RECT 121.385 207.275 121.765 207.655 ;
        RECT 123.235 207.155 123.550 211.480 ;
        RECT 123.845 209.230 124.125 210.760 ;
        RECT 124.415 205.915 124.715 212.955 ;
        RECT 126.190 206.670 126.490 210.730 ;
        RECT 123.710 204.105 124.090 204.485 ;
        RECT 127.440 203.700 127.730 212.945 ;
        RECT 129.290 205.400 129.590 212.210 ;
        RECT 130.080 205.995 130.390 214.730 ;
        RECT 130.875 205.925 131.175 212.755 ;
        RECT 132.680 206.655 132.960 210.745 ;
        RECT 133.450 205.185 133.730 208.220 ;
        RECT 136.200 205.140 136.500 212.295 ;
        RECT 138.540 210.910 138.915 219.110 ;
        RECT 140.285 210.105 140.585 221.100 ;
        RECT 11.820 185.655 12.120 192.585 ;
        RECT 13.130 186.255 13.430 192.605 ;
        RECT 14.445 186.285 14.740 193.110 ;
        RECT 18.285 185.655 18.585 192.595 ;
        RECT 20.495 186.230 20.800 192.590 ;
        RECT 21.345 186.230 21.645 193.050 ;
        RECT 23.155 189.675 23.535 190.055 ;
        RECT 24.940 188.255 25.260 190.385 ;
        RECT 23.370 184.965 23.750 187.985 ;
        RECT 25.550 187.415 25.830 189.820 ;
        RECT 26.160 186.260 26.460 193.300 ;
        RECT 27.280 185.655 27.580 192.585 ;
        RECT 28.590 186.255 28.890 192.605 ;
        RECT 29.185 188.130 29.510 193.290 ;
        RECT 29.905 186.285 30.200 193.110 ;
        RECT 31.035 185.745 31.335 192.555 ;
        RECT 31.825 186.340 32.135 192.530 ;
        RECT 32.620 186.270 32.920 193.100 ;
        RECT 33.745 185.655 34.045 192.595 ;
        RECT 35.195 185.530 35.475 188.565 ;
        RECT 35.955 186.230 36.275 192.590 ;
        RECT 36.805 186.230 37.105 193.050 ;
        RECT 37.945 185.485 38.245 192.640 ;
        RECT 38.580 187.630 38.960 188.010 ;
        RECT 39.285 183.515 39.645 190.075 ;
        RECT 40.425 188.265 40.750 190.130 ;
        RECT 41.090 184.920 41.550 189.605 ;
        RECT 41.875 187.465 42.325 196.285 ;
        RECT 44.060 189.290 44.490 192.280 ;
        RECT 41.805 183.575 42.185 183.955 ;
        RECT 44.695 183.595 45.075 184.970 ;
        RECT 45.465 184.415 45.780 195.465 ;
        RECT 46.480 194.160 46.770 196.220 ;
        RECT 46.400 186.305 46.725 188.675 ;
        RECT 48.050 188.350 48.450 192.315 ;
        RECT 48.770 184.245 49.095 187.010 ;
        RECT 49.755 186.280 50.160 189.610 ;
        RECT 54.405 183.305 54.775 192.405 ;
        RECT 55.350 184.370 55.640 196.205 ;
        RECT 63.255 194.100 63.565 196.615 ;
        RECT 59.165 186.335 59.605 189.610 ;
        RECT 61.545 188.350 62.070 192.290 ;
        RECT 60.705 184.245 61.030 187.010 ;
        RECT 63.220 186.340 63.635 188.730 ;
        RECT 64.250 184.900 64.565 195.585 ;
        RECT 65.580 189.290 66.065 192.300 ;
        RECT 64.950 183.510 65.285 184.860 ;
        RECT 5.160 167.355 5.575 181.080 ;
        RECT 68.475 180.300 69.030 191.315 ;
        RECT 6.600 168.380 7.015 179.745 ;
        RECT 69.705 178.895 70.175 188.240 ;
        RECT 75.485 179.070 76.010 190.490 ;
        RECT 77.615 180.475 78.080 191.815 ;
        RECT 81.435 184.425 81.790 195.510 ;
        RECT 85.180 194.150 85.470 196.210 ;
        RECT 91.960 193.000 92.270 193.030 ;
        RECT 82.760 189.280 83.230 192.270 ;
        RECT 85.110 186.295 85.425 188.665 ;
        RECT 86.730 188.340 87.150 192.305 ;
        RECT 83.395 183.585 83.775 184.960 ;
        RECT 87.470 184.235 87.795 187.000 ;
        RECT 88.455 186.270 88.860 189.600 ;
        RECT 91.960 186.900 92.275 193.000 ;
        RECT 93.105 183.295 93.475 192.395 ;
        RECT 94.050 184.360 94.340 196.195 ;
        RECT 101.955 194.090 102.265 196.605 ;
        RECT 106.205 195.790 106.585 196.170 ;
        RECT 108.335 195.790 108.715 196.170 ;
        RECT 94.945 186.855 95.275 193.050 ;
        RECT 97.850 186.325 98.305 189.600 ;
        RECT 100.210 188.340 100.755 192.280 ;
        RECT 104.265 189.280 104.700 192.290 ;
        RECT 99.405 184.235 99.730 187.000 ;
        RECT 101.920 186.330 102.335 188.720 ;
        RECT 105.460 184.905 105.790 195.600 ;
        RECT 106.895 189.240 107.280 195.025 ;
        RECT 103.650 183.500 103.985 184.850 ;
        RECT 107.255 184.485 107.680 188.760 ;
        RECT 108.955 186.250 109.255 193.290 ;
        RECT 110.075 185.645 110.375 192.575 ;
        RECT 111.385 186.245 111.685 192.595 ;
        RECT 105.915 183.575 106.295 183.955 ;
        RECT 108.110 183.560 108.490 183.940 ;
        RECT 111.980 183.500 112.270 193.280 ;
        RECT 112.700 186.275 112.995 193.100 ;
        RECT 113.830 185.735 114.130 192.545 ;
        RECT 114.620 186.330 114.930 196.370 ;
        RECT 123.810 194.615 124.190 194.995 ;
        RECT 115.415 186.260 115.715 193.090 ;
        RECT 116.540 185.645 116.840 192.585 ;
        RECT 117.990 185.520 118.270 188.555 ;
        RECT 118.750 186.220 119.030 192.580 ;
        RECT 119.600 186.220 119.900 193.040 ;
        RECT 120.740 185.475 121.040 192.630 ;
        RECT 121.385 189.665 121.765 190.045 ;
        RECT 121.385 187.610 121.765 187.990 ;
        RECT 123.235 187.490 123.550 191.815 ;
        RECT 123.845 189.565 124.125 191.095 ;
        RECT 124.415 186.250 124.715 193.290 ;
        RECT 126.190 187.005 126.490 191.065 ;
        RECT 123.710 184.440 124.090 184.820 ;
        RECT 127.440 184.035 127.730 193.280 ;
        RECT 129.290 185.735 129.590 192.545 ;
        RECT 130.080 186.330 130.390 195.065 ;
        RECT 130.875 186.260 131.175 193.090 ;
        RECT 132.680 186.990 132.960 191.080 ;
        RECT 133.450 185.520 133.730 188.555 ;
        RECT 136.200 185.475 136.500 192.630 ;
        RECT 138.125 191.395 138.500 199.235 ;
        RECT 139.980 190.645 140.280 201.185 ;
        RECT 11.970 165.860 12.270 172.790 ;
        RECT 13.280 166.460 13.580 172.810 ;
        RECT 14.595 166.490 14.890 173.315 ;
        RECT 18.435 165.860 18.735 172.800 ;
        RECT 20.645 166.435 20.950 172.795 ;
        RECT 21.495 166.435 21.795 173.255 ;
        RECT 23.305 169.880 23.685 170.260 ;
        RECT 25.090 168.460 25.410 170.590 ;
        RECT 23.520 165.170 23.900 168.190 ;
        RECT 25.700 167.620 25.980 170.025 ;
        RECT 26.310 166.465 26.610 173.505 ;
        RECT 27.430 165.860 27.730 172.790 ;
        RECT 28.740 166.460 29.040 172.810 ;
        RECT 29.335 168.335 29.660 173.495 ;
        RECT 30.055 166.490 30.350 173.315 ;
        RECT 31.185 165.950 31.485 172.760 ;
        RECT 31.975 166.545 32.285 172.735 ;
        RECT 32.770 166.475 33.070 173.305 ;
        RECT 33.895 165.860 34.195 172.800 ;
        RECT 35.345 165.735 35.625 168.770 ;
        RECT 36.105 166.435 36.425 172.795 ;
        RECT 36.955 166.435 37.255 173.255 ;
        RECT 38.095 165.690 38.395 172.845 ;
        RECT 38.730 167.835 39.110 168.215 ;
        RECT 39.435 163.720 39.795 170.280 ;
        RECT 40.575 168.470 40.900 170.335 ;
        RECT 41.240 165.125 41.700 169.810 ;
        RECT 42.025 167.670 42.475 176.490 ;
        RECT 44.210 169.495 44.640 172.485 ;
        RECT 41.955 163.780 42.335 164.160 ;
        RECT 44.845 163.800 45.225 165.175 ;
        RECT 45.615 164.620 45.930 175.670 ;
        RECT 46.630 174.365 46.920 176.425 ;
        RECT 46.550 166.510 46.875 168.880 ;
        RECT 48.200 168.555 48.600 172.520 ;
        RECT 48.920 164.450 49.245 167.215 ;
        RECT 49.905 166.485 50.310 169.815 ;
        RECT 54.555 163.510 54.925 172.610 ;
        RECT 55.500 164.575 55.790 176.410 ;
        RECT 63.405 174.305 63.715 176.820 ;
        RECT 59.315 166.540 59.755 169.815 ;
        RECT 61.695 168.555 62.220 172.495 ;
        RECT 60.855 164.450 61.180 167.215 ;
        RECT 63.370 166.545 63.785 168.935 ;
        RECT 64.400 165.105 64.715 175.790 ;
        RECT 65.730 169.495 66.215 172.505 ;
        RECT 65.100 163.715 65.435 165.065 ;
        RECT 4.815 147.890 5.170 161.680 ;
        RECT 68.160 161.050 68.610 171.315 ;
        RECT 6.440 148.745 6.800 160.080 ;
        RECT 69.325 159.510 69.810 168.395 ;
        RECT 75.630 159.135 76.035 170.665 ;
        RECT 77.705 161.035 78.095 172.135 ;
        RECT 81.475 164.585 81.830 175.670 ;
        RECT 85.220 174.310 85.510 176.370 ;
        RECT 92.000 173.160 92.310 173.190 ;
        RECT 82.800 169.440 83.270 172.430 ;
        RECT 85.150 166.455 85.465 168.825 ;
        RECT 86.770 168.500 87.190 172.465 ;
        RECT 83.435 163.745 83.815 165.120 ;
        RECT 87.510 164.395 87.835 167.160 ;
        RECT 88.495 166.430 88.900 169.760 ;
        RECT 92.000 167.060 92.315 173.160 ;
        RECT 93.145 163.455 93.515 172.555 ;
        RECT 94.090 164.520 94.380 176.355 ;
        RECT 101.995 174.250 102.305 176.765 ;
        RECT 106.245 175.950 106.625 176.330 ;
        RECT 108.375 175.950 108.755 176.330 ;
        RECT 94.985 167.015 95.315 173.210 ;
        RECT 97.890 166.485 98.345 169.760 ;
        RECT 100.250 168.500 100.795 172.440 ;
        RECT 104.305 169.440 104.740 172.450 ;
        RECT 99.445 164.395 99.770 167.160 ;
        RECT 101.960 166.490 102.375 168.880 ;
        RECT 105.500 165.065 105.830 175.760 ;
        RECT 106.935 169.400 107.320 175.185 ;
        RECT 103.690 163.660 104.025 165.010 ;
        RECT 107.295 164.645 107.720 168.920 ;
        RECT 108.995 166.410 109.295 173.450 ;
        RECT 110.115 165.805 110.415 172.735 ;
        RECT 111.425 166.405 111.725 172.755 ;
        RECT 105.955 163.735 106.335 164.115 ;
        RECT 108.150 163.720 108.530 164.100 ;
        RECT 112.020 163.660 112.310 173.440 ;
        RECT 112.740 166.435 113.035 173.260 ;
        RECT 113.870 165.895 114.170 172.705 ;
        RECT 114.660 166.490 114.970 176.530 ;
        RECT 123.850 174.775 124.230 175.155 ;
        RECT 115.455 166.420 115.755 173.250 ;
        RECT 116.580 165.805 116.880 172.745 ;
        RECT 118.030 165.680 118.310 168.715 ;
        RECT 118.790 166.380 119.070 172.740 ;
        RECT 119.640 166.380 119.940 173.200 ;
        RECT 120.780 165.635 121.080 172.790 ;
        RECT 121.425 169.825 121.805 170.205 ;
        RECT 121.425 167.770 121.805 168.150 ;
        RECT 123.275 167.650 123.590 171.975 ;
        RECT 123.885 169.725 124.165 171.255 ;
        RECT 124.455 166.410 124.755 173.450 ;
        RECT 126.230 167.165 126.530 171.225 ;
        RECT 123.750 164.600 124.130 164.980 ;
        RECT 127.480 164.195 127.770 173.440 ;
        RECT 129.330 165.895 129.630 172.705 ;
        RECT 130.120 166.490 130.430 175.225 ;
        RECT 130.915 166.420 131.215 173.250 ;
        RECT 132.720 167.150 133.000 171.240 ;
        RECT 133.490 165.680 133.770 168.715 ;
        RECT 136.240 165.635 136.540 172.790 ;
        RECT 138.440 171.420 138.840 180.160 ;
        RECT 140.020 170.640 140.415 181.520 ;
        RECT 11.925 146.170 12.225 153.100 ;
        RECT 13.235 146.770 13.535 153.120 ;
        RECT 14.550 146.800 14.845 153.625 ;
        RECT 18.390 146.170 18.690 153.110 ;
        RECT 20.600 146.745 20.905 153.105 ;
        RECT 21.450 146.745 21.750 153.565 ;
        RECT 23.260 150.190 23.640 150.570 ;
        RECT 25.045 148.770 25.365 150.900 ;
        RECT 23.475 145.480 23.855 148.500 ;
        RECT 25.655 147.930 25.935 150.335 ;
        RECT 26.265 146.775 26.565 153.815 ;
        RECT 27.385 146.170 27.685 153.100 ;
        RECT 28.695 146.770 28.995 153.120 ;
        RECT 29.290 148.645 29.615 153.805 ;
        RECT 30.010 146.800 30.305 153.625 ;
        RECT 31.140 146.260 31.440 153.070 ;
        RECT 31.930 146.855 32.240 153.045 ;
        RECT 32.725 146.785 33.025 153.615 ;
        RECT 33.850 146.170 34.150 153.110 ;
        RECT 35.300 146.045 35.580 149.080 ;
        RECT 36.060 146.745 36.380 153.105 ;
        RECT 36.910 146.745 37.210 153.565 ;
        RECT 38.050 146.000 38.350 153.155 ;
        RECT 38.685 148.145 39.065 148.525 ;
        RECT 39.390 144.030 39.750 150.590 ;
        RECT 40.530 148.780 40.855 150.645 ;
        RECT 41.195 145.435 41.655 150.120 ;
        RECT 41.980 147.980 42.430 156.800 ;
        RECT 44.165 149.805 44.595 152.795 ;
        RECT 41.910 144.090 42.290 144.470 ;
        RECT 44.800 144.110 45.180 145.485 ;
        RECT 45.570 144.930 45.885 155.980 ;
        RECT 46.585 154.675 46.875 156.735 ;
        RECT 46.505 146.820 46.830 149.190 ;
        RECT 48.155 148.865 48.555 152.830 ;
        RECT 48.875 144.760 49.200 147.525 ;
        RECT 49.860 146.795 50.265 150.125 ;
        RECT 54.510 143.820 54.880 152.920 ;
        RECT 55.455 144.885 55.745 156.720 ;
        RECT 63.360 154.615 63.670 157.130 ;
        RECT 59.270 146.850 59.710 150.125 ;
        RECT 61.650 148.865 62.175 152.805 ;
        RECT 60.810 144.760 61.135 147.525 ;
        RECT 63.325 146.855 63.740 149.245 ;
        RECT 64.355 145.415 64.670 156.100 ;
        RECT 65.685 149.805 66.170 152.815 ;
        RECT 65.055 144.025 65.390 145.375 ;
        RECT 4.815 128.125 5.170 142.180 ;
        RECT 68.160 141.550 68.610 151.665 ;
        RECT 6.440 128.930 6.800 140.580 ;
        RECT 69.325 140.010 69.810 148.765 ;
        RECT 75.930 139.385 76.335 150.915 ;
        RECT 78.005 141.285 78.395 152.385 ;
        RECT 81.275 144.860 81.630 155.945 ;
        RECT 85.020 154.585 85.310 156.645 ;
        RECT 91.800 153.435 92.110 153.465 ;
        RECT 82.600 149.715 83.070 152.705 ;
        RECT 84.950 146.730 85.265 149.100 ;
        RECT 86.570 148.775 86.990 152.740 ;
        RECT 83.235 144.020 83.615 145.395 ;
        RECT 87.310 144.670 87.635 147.435 ;
        RECT 88.295 146.705 88.700 150.035 ;
        RECT 91.800 147.335 92.115 153.435 ;
        RECT 92.945 143.730 93.315 152.830 ;
        RECT 93.890 144.795 94.180 156.630 ;
        RECT 101.795 154.525 102.105 157.040 ;
        RECT 106.045 156.225 106.425 156.605 ;
        RECT 108.175 156.225 108.555 156.605 ;
        RECT 94.785 147.290 95.115 153.485 ;
        RECT 97.690 146.760 98.145 150.035 ;
        RECT 100.050 148.775 100.595 152.715 ;
        RECT 104.105 149.715 104.540 152.725 ;
        RECT 99.245 144.670 99.570 147.435 ;
        RECT 101.760 146.765 102.175 149.155 ;
        RECT 105.300 145.340 105.630 156.035 ;
        RECT 106.735 149.675 107.120 155.460 ;
        RECT 103.490 143.935 103.825 145.285 ;
        RECT 107.095 144.920 107.520 149.195 ;
        RECT 108.795 146.685 109.095 153.725 ;
        RECT 109.915 146.080 110.215 153.010 ;
        RECT 111.225 146.680 111.525 153.030 ;
        RECT 105.755 144.010 106.135 144.390 ;
        RECT 107.950 143.995 108.330 144.375 ;
        RECT 111.820 143.935 112.110 153.715 ;
        RECT 112.540 146.710 112.835 153.535 ;
        RECT 113.670 146.170 113.970 152.980 ;
        RECT 114.460 146.765 114.770 156.805 ;
        RECT 123.650 155.050 124.030 155.430 ;
        RECT 115.255 146.695 115.555 153.525 ;
        RECT 116.380 146.080 116.680 153.020 ;
        RECT 117.830 145.955 118.110 148.990 ;
        RECT 118.590 146.655 118.870 153.015 ;
        RECT 119.440 146.655 119.740 153.475 ;
        RECT 120.580 145.910 120.880 153.065 ;
        RECT 121.225 150.100 121.605 150.480 ;
        RECT 121.225 148.045 121.605 148.425 ;
        RECT 123.075 147.925 123.390 152.250 ;
        RECT 123.685 150.000 123.965 151.530 ;
        RECT 124.255 146.685 124.555 153.725 ;
        RECT 126.030 147.440 126.330 151.500 ;
        RECT 123.550 144.875 123.930 145.255 ;
        RECT 127.280 144.470 127.570 153.715 ;
        RECT 129.130 146.170 129.430 152.980 ;
        RECT 129.920 146.765 130.230 155.500 ;
        RECT 130.715 146.695 131.015 153.525 ;
        RECT 132.520 147.425 132.800 151.515 ;
        RECT 133.290 145.955 133.570 148.990 ;
        RECT 136.040 145.910 136.340 153.065 ;
        RECT 138.080 151.805 138.455 160.005 ;
        RECT 139.825 151.000 140.125 161.995 ;
        RECT 12.115 126.460 12.415 133.390 ;
        RECT 13.425 127.060 13.725 133.410 ;
        RECT 14.740 127.090 15.035 133.915 ;
        RECT 18.580 126.460 18.880 133.400 ;
        RECT 20.790 127.035 21.095 133.395 ;
        RECT 21.640 127.035 21.940 133.855 ;
        RECT 23.450 130.480 23.830 130.860 ;
        RECT 25.235 129.060 25.555 131.190 ;
        RECT 23.665 125.770 24.045 128.790 ;
        RECT 25.845 128.220 26.125 130.625 ;
        RECT 26.455 127.065 26.755 134.105 ;
        RECT 27.575 126.460 27.875 133.390 ;
        RECT 28.885 127.060 29.185 133.410 ;
        RECT 29.480 128.935 29.805 134.095 ;
        RECT 30.200 127.090 30.495 133.915 ;
        RECT 31.330 126.550 31.630 133.360 ;
        RECT 32.120 127.145 32.430 133.335 ;
        RECT 32.915 127.075 33.215 133.905 ;
        RECT 34.040 126.460 34.340 133.400 ;
        RECT 35.490 126.335 35.770 129.370 ;
        RECT 36.250 127.035 36.570 133.395 ;
        RECT 37.100 127.035 37.400 133.855 ;
        RECT 38.240 126.290 38.540 133.445 ;
        RECT 38.875 128.435 39.255 128.815 ;
        RECT 39.580 124.320 39.940 130.880 ;
        RECT 40.720 129.070 41.045 130.935 ;
        RECT 41.385 125.725 41.845 130.410 ;
        RECT 42.170 128.270 42.620 137.090 ;
        RECT 44.355 130.095 44.785 133.085 ;
        RECT 42.100 124.380 42.480 124.760 ;
        RECT 44.990 124.400 45.370 125.775 ;
        RECT 45.760 125.220 46.075 136.270 ;
        RECT 46.775 134.965 47.065 137.025 ;
        RECT 46.695 127.110 47.020 129.480 ;
        RECT 48.345 129.155 48.745 133.120 ;
        RECT 49.065 125.050 49.390 127.815 ;
        RECT 50.050 127.085 50.455 130.415 ;
        RECT 54.700 124.110 55.070 133.210 ;
        RECT 55.645 125.175 55.935 137.010 ;
        RECT 63.550 134.905 63.860 137.420 ;
        RECT 59.460 127.140 59.900 130.415 ;
        RECT 61.840 129.155 62.365 133.095 ;
        RECT 61.000 125.050 61.325 127.815 ;
        RECT 63.515 127.145 63.930 129.535 ;
        RECT 64.545 125.705 64.860 136.390 ;
        RECT 65.875 130.095 66.360 133.105 ;
        RECT 65.245 124.315 65.580 125.665 ;
        RECT 5.025 108.350 5.380 122.140 ;
        RECT 68.370 121.510 68.820 132.010 ;
        RECT 6.650 109.205 7.010 120.540 ;
        RECT 69.535 119.970 70.020 129.210 ;
        RECT 75.950 119.725 76.355 131.255 ;
        RECT 78.025 121.625 78.415 132.725 ;
        RECT 81.430 125.215 81.785 136.300 ;
        RECT 85.175 134.940 85.465 137.000 ;
        RECT 91.955 133.790 92.265 133.820 ;
        RECT 82.755 130.070 83.225 133.060 ;
        RECT 85.105 127.085 85.420 129.455 ;
        RECT 86.725 129.130 87.145 133.095 ;
        RECT 83.390 124.375 83.770 125.750 ;
        RECT 87.465 125.025 87.790 127.790 ;
        RECT 88.450 127.060 88.855 130.390 ;
        RECT 91.955 127.690 92.270 133.790 ;
        RECT 93.100 124.085 93.470 133.185 ;
        RECT 94.045 125.150 94.335 136.985 ;
        RECT 101.950 134.880 102.260 137.395 ;
        RECT 106.200 136.580 106.580 136.960 ;
        RECT 108.330 136.580 108.710 136.960 ;
        RECT 94.940 127.645 95.270 133.840 ;
        RECT 97.845 127.115 98.300 130.390 ;
        RECT 100.205 129.130 100.750 133.070 ;
        RECT 104.260 130.070 104.695 133.080 ;
        RECT 99.400 125.025 99.725 127.790 ;
        RECT 101.915 127.120 102.330 129.510 ;
        RECT 105.455 125.695 105.785 136.390 ;
        RECT 106.890 130.030 107.275 135.815 ;
        RECT 103.645 124.290 103.980 125.640 ;
        RECT 107.250 125.275 107.675 129.550 ;
        RECT 108.950 127.040 109.250 134.080 ;
        RECT 110.070 126.435 110.370 133.365 ;
        RECT 111.380 127.035 111.680 133.385 ;
        RECT 105.910 124.365 106.290 124.745 ;
        RECT 108.105 124.350 108.485 124.730 ;
        RECT 111.975 124.290 112.265 134.070 ;
        RECT 112.695 127.065 112.990 133.890 ;
        RECT 113.825 126.525 114.125 133.335 ;
        RECT 114.615 127.120 114.925 137.160 ;
        RECT 123.805 135.405 124.185 135.785 ;
        RECT 115.410 127.050 115.710 133.880 ;
        RECT 116.535 126.435 116.835 133.375 ;
        RECT 117.985 126.310 118.265 129.345 ;
        RECT 118.745 127.010 119.025 133.370 ;
        RECT 119.595 127.010 119.895 133.830 ;
        RECT 120.735 126.265 121.035 133.420 ;
        RECT 121.380 130.455 121.760 130.835 ;
        RECT 121.380 128.400 121.760 128.780 ;
        RECT 123.230 128.280 123.545 132.605 ;
        RECT 123.840 130.355 124.120 131.885 ;
        RECT 124.410 127.040 124.710 134.080 ;
        RECT 126.185 127.795 126.485 131.855 ;
        RECT 123.705 125.230 124.085 125.610 ;
        RECT 127.435 124.825 127.725 134.070 ;
        RECT 129.285 126.525 129.585 133.335 ;
        RECT 130.075 127.120 130.385 135.855 ;
        RECT 130.870 127.050 131.170 133.880 ;
        RECT 132.675 127.780 132.955 131.870 ;
        RECT 133.445 126.310 133.725 129.345 ;
        RECT 136.195 126.265 136.495 133.420 ;
        RECT 138.380 132.055 138.755 140.255 ;
        RECT 140.125 131.250 140.425 142.245 ;
        RECT 11.920 106.620 12.220 113.550 ;
        RECT 13.230 107.220 13.530 113.570 ;
        RECT 14.545 107.250 14.840 114.075 ;
        RECT 18.385 106.620 18.685 113.560 ;
        RECT 20.595 107.195 20.900 113.555 ;
        RECT 21.445 107.195 21.745 114.015 ;
        RECT 23.255 110.640 23.635 111.020 ;
        RECT 25.040 109.220 25.360 111.350 ;
        RECT 23.470 105.930 23.850 108.950 ;
        RECT 25.650 108.380 25.930 110.785 ;
        RECT 26.260 107.225 26.560 114.265 ;
        RECT 27.380 106.620 27.680 113.550 ;
        RECT 28.690 107.220 28.990 113.570 ;
        RECT 29.285 109.095 29.610 114.255 ;
        RECT 30.005 107.250 30.300 114.075 ;
        RECT 31.135 106.710 31.435 113.520 ;
        RECT 31.925 107.305 32.235 113.495 ;
        RECT 32.720 107.235 33.020 114.065 ;
        RECT 33.845 106.620 34.145 113.560 ;
        RECT 35.295 106.495 35.575 109.530 ;
        RECT 36.055 107.195 36.375 113.555 ;
        RECT 36.905 107.195 37.205 114.015 ;
        RECT 38.045 106.450 38.345 113.605 ;
        RECT 38.680 108.595 39.060 108.975 ;
        RECT 39.385 104.480 39.745 111.040 ;
        RECT 40.525 109.230 40.850 111.095 ;
        RECT 41.190 105.885 41.650 110.570 ;
        RECT 41.975 108.430 42.425 117.250 ;
        RECT 44.160 110.255 44.590 113.245 ;
        RECT 41.905 104.540 42.285 104.920 ;
        RECT 44.795 104.560 45.175 105.935 ;
        RECT 45.565 105.380 45.880 116.430 ;
        RECT 46.580 115.125 46.870 117.185 ;
        RECT 46.500 107.270 46.825 109.640 ;
        RECT 48.150 109.315 48.550 113.280 ;
        RECT 48.870 105.210 49.195 107.975 ;
        RECT 49.855 107.245 50.260 110.575 ;
        RECT 54.505 104.270 54.875 113.370 ;
        RECT 55.450 105.335 55.740 117.170 ;
        RECT 63.355 115.065 63.665 117.580 ;
        RECT 59.265 107.300 59.705 110.575 ;
        RECT 61.645 109.315 62.170 113.255 ;
        RECT 60.805 105.210 61.130 107.975 ;
        RECT 63.320 107.305 63.735 109.695 ;
        RECT 64.350 105.865 64.665 116.550 ;
        RECT 65.680 110.255 66.165 113.265 ;
        RECT 65.050 104.475 65.385 105.825 ;
        RECT 4.980 88.560 5.335 102.350 ;
        RECT 68.325 101.720 68.775 112.210 ;
        RECT 6.605 89.465 6.965 100.750 ;
        RECT 69.490 100.180 69.975 109.340 ;
        RECT 75.950 99.990 76.355 111.520 ;
        RECT 78.025 101.890 78.415 112.990 ;
        RECT 81.430 105.420 81.785 116.505 ;
        RECT 85.175 115.145 85.465 117.205 ;
        RECT 91.955 113.995 92.265 114.025 ;
        RECT 82.755 110.275 83.225 113.265 ;
        RECT 85.105 107.290 85.420 109.660 ;
        RECT 86.725 109.335 87.145 113.300 ;
        RECT 83.390 104.580 83.770 105.955 ;
        RECT 87.465 105.230 87.790 107.995 ;
        RECT 88.450 107.265 88.855 110.595 ;
        RECT 91.955 107.895 92.270 113.995 ;
        RECT 93.100 104.290 93.470 113.390 ;
        RECT 94.045 105.355 94.335 117.190 ;
        RECT 101.950 115.085 102.260 117.600 ;
        RECT 106.200 116.785 106.580 117.165 ;
        RECT 108.330 116.785 108.710 117.165 ;
        RECT 94.940 107.850 95.270 114.045 ;
        RECT 97.845 107.320 98.300 110.595 ;
        RECT 100.205 109.335 100.750 113.275 ;
        RECT 104.260 110.275 104.695 113.285 ;
        RECT 99.400 105.230 99.725 107.995 ;
        RECT 101.915 107.325 102.330 109.715 ;
        RECT 105.455 105.900 105.785 116.595 ;
        RECT 106.890 110.235 107.275 116.020 ;
        RECT 103.645 104.495 103.980 105.845 ;
        RECT 107.250 105.480 107.675 109.755 ;
        RECT 108.950 107.245 109.250 114.285 ;
        RECT 110.070 106.640 110.370 113.570 ;
        RECT 111.380 107.240 111.680 113.590 ;
        RECT 105.910 104.570 106.290 104.950 ;
        RECT 108.105 104.555 108.485 104.935 ;
        RECT 111.975 104.495 112.265 114.275 ;
        RECT 112.695 107.270 112.990 114.095 ;
        RECT 113.825 106.730 114.125 113.540 ;
        RECT 114.615 107.325 114.925 117.365 ;
        RECT 123.805 115.610 124.185 115.990 ;
        RECT 115.410 107.255 115.710 114.085 ;
        RECT 116.535 106.640 116.835 113.580 ;
        RECT 117.985 106.515 118.265 109.550 ;
        RECT 118.745 107.215 119.025 113.575 ;
        RECT 119.595 107.215 119.895 114.035 ;
        RECT 120.735 106.470 121.035 113.625 ;
        RECT 121.380 110.660 121.760 111.040 ;
        RECT 121.380 108.605 121.760 108.985 ;
        RECT 123.230 108.485 123.545 112.810 ;
        RECT 123.840 110.560 124.120 112.090 ;
        RECT 124.410 107.245 124.710 114.285 ;
        RECT 126.185 108.000 126.485 112.060 ;
        RECT 123.705 105.435 124.085 105.815 ;
        RECT 127.435 105.030 127.725 114.275 ;
        RECT 129.285 106.730 129.585 113.540 ;
        RECT 130.075 107.325 130.385 116.060 ;
        RECT 130.870 107.255 131.170 114.085 ;
        RECT 132.675 107.985 132.955 112.075 ;
        RECT 133.445 106.515 133.725 109.550 ;
        RECT 136.195 106.470 136.495 113.625 ;
        RECT 138.400 112.395 138.775 120.595 ;
        RECT 140.145 111.590 140.445 122.585 ;
        RECT 11.790 86.910 12.090 93.840 ;
        RECT 13.100 87.510 13.400 93.860 ;
        RECT 14.415 87.540 14.710 94.365 ;
        RECT 18.255 86.910 18.555 93.850 ;
        RECT 20.465 87.485 20.770 93.845 ;
        RECT 21.315 87.485 21.615 94.305 ;
        RECT 23.125 90.930 23.505 91.310 ;
        RECT 24.910 89.510 25.230 91.640 ;
        RECT 23.340 86.220 23.720 89.240 ;
        RECT 25.520 88.670 25.800 91.075 ;
        RECT 26.130 87.515 26.430 94.555 ;
        RECT 27.250 86.910 27.550 93.840 ;
        RECT 28.560 87.510 28.860 93.860 ;
        RECT 29.155 89.385 29.480 94.545 ;
        RECT 29.875 87.540 30.170 94.365 ;
        RECT 31.005 87.000 31.305 93.810 ;
        RECT 31.795 87.595 32.105 93.785 ;
        RECT 32.590 87.525 32.890 94.355 ;
        RECT 33.715 86.910 34.015 93.850 ;
        RECT 35.165 86.785 35.445 89.820 ;
        RECT 35.925 87.485 36.245 93.845 ;
        RECT 36.775 87.485 37.075 94.305 ;
        RECT 37.915 86.740 38.215 93.895 ;
        RECT 38.550 88.885 38.930 89.265 ;
        RECT 39.255 84.770 39.615 91.330 ;
        RECT 40.395 89.520 40.720 91.385 ;
        RECT 41.060 86.175 41.520 90.860 ;
        RECT 41.845 88.720 42.295 97.540 ;
        RECT 44.030 90.545 44.460 93.535 ;
        RECT 41.775 84.830 42.155 85.210 ;
        RECT 44.665 84.850 45.045 86.225 ;
        RECT 45.435 85.670 45.750 96.720 ;
        RECT 46.450 95.415 46.740 97.475 ;
        RECT 46.370 87.560 46.695 89.930 ;
        RECT 48.020 89.605 48.420 93.570 ;
        RECT 48.740 85.500 49.065 88.265 ;
        RECT 49.725 87.535 50.130 90.865 ;
        RECT 54.375 84.560 54.745 93.660 ;
        RECT 55.320 85.625 55.610 97.460 ;
        RECT 63.225 95.355 63.535 97.870 ;
        RECT 59.135 87.590 59.575 90.865 ;
        RECT 61.515 89.605 62.040 93.545 ;
        RECT 60.675 85.500 61.000 88.265 ;
        RECT 63.190 87.595 63.605 89.985 ;
        RECT 64.220 86.155 64.535 96.840 ;
        RECT 65.550 90.545 66.035 93.555 ;
        RECT 64.920 84.765 65.255 86.115 ;
        RECT 4.675 68.800 5.030 82.720 ;
        RECT 68.020 82.090 68.470 92.355 ;
        RECT 6.300 69.705 6.660 81.120 ;
        RECT 69.185 80.550 69.670 89.435 ;
        RECT 75.850 80.285 76.255 91.815 ;
        RECT 77.925 82.185 78.315 93.285 ;
        RECT 81.350 85.665 81.705 96.750 ;
        RECT 85.095 95.390 85.385 97.450 ;
        RECT 91.875 94.240 92.185 94.270 ;
        RECT 82.675 90.520 83.145 93.510 ;
        RECT 85.025 87.535 85.340 89.905 ;
        RECT 86.645 89.580 87.065 93.545 ;
        RECT 83.310 84.825 83.690 86.200 ;
        RECT 87.385 85.475 87.710 88.240 ;
        RECT 88.370 87.510 88.775 90.840 ;
        RECT 91.875 88.140 92.190 94.240 ;
        RECT 93.020 84.535 93.390 93.635 ;
        RECT 93.965 85.600 94.255 97.435 ;
        RECT 101.870 95.330 102.180 97.845 ;
        RECT 106.120 97.030 106.500 97.410 ;
        RECT 108.250 97.030 108.630 97.410 ;
        RECT 94.860 88.095 95.190 94.290 ;
        RECT 97.765 87.565 98.220 90.840 ;
        RECT 100.125 89.580 100.670 93.520 ;
        RECT 104.180 90.520 104.615 93.530 ;
        RECT 99.320 85.475 99.645 88.240 ;
        RECT 101.835 87.570 102.250 89.960 ;
        RECT 105.375 86.145 105.705 96.840 ;
        RECT 106.810 90.480 107.195 96.265 ;
        RECT 103.565 84.740 103.900 86.090 ;
        RECT 107.170 85.725 107.595 90.000 ;
        RECT 108.870 87.490 109.170 94.530 ;
        RECT 109.990 86.885 110.290 93.815 ;
        RECT 111.300 87.485 111.600 93.835 ;
        RECT 105.830 84.815 106.210 85.195 ;
        RECT 108.025 84.800 108.405 85.180 ;
        RECT 111.895 84.740 112.185 94.520 ;
        RECT 112.615 87.515 112.910 94.340 ;
        RECT 113.745 86.975 114.045 93.785 ;
        RECT 114.535 87.570 114.845 97.610 ;
        RECT 123.725 95.855 124.105 96.235 ;
        RECT 115.330 87.500 115.630 94.330 ;
        RECT 116.455 86.885 116.755 93.825 ;
        RECT 117.905 86.760 118.185 89.795 ;
        RECT 118.665 87.460 118.945 93.820 ;
        RECT 119.515 87.460 119.815 94.280 ;
        RECT 120.655 86.715 120.955 93.870 ;
        RECT 121.300 90.905 121.680 91.285 ;
        RECT 121.300 88.850 121.680 89.230 ;
        RECT 123.150 88.730 123.465 93.055 ;
        RECT 123.760 90.805 124.040 92.335 ;
        RECT 124.330 87.490 124.630 94.530 ;
        RECT 126.105 88.245 126.405 92.305 ;
        RECT 123.625 85.680 124.005 86.060 ;
        RECT 127.355 85.275 127.645 94.520 ;
        RECT 129.205 86.975 129.505 93.785 ;
        RECT 129.995 87.570 130.305 96.305 ;
        RECT 130.790 87.500 131.090 94.330 ;
        RECT 132.595 88.230 132.875 92.320 ;
        RECT 133.365 86.760 133.645 89.795 ;
        RECT 136.115 86.715 136.415 93.870 ;
        RECT 138.400 92.575 138.775 100.860 ;
        RECT 140.145 91.855 140.445 102.850 ;
        RECT 11.920 67.150 12.220 74.080 ;
        RECT 13.230 67.750 13.530 74.100 ;
        RECT 14.545 67.780 14.840 74.605 ;
        RECT 18.385 67.150 18.685 74.090 ;
        RECT 20.595 67.725 20.900 74.085 ;
        RECT 21.445 67.725 21.745 74.545 ;
        RECT 23.255 71.170 23.635 71.550 ;
        RECT 25.040 69.750 25.360 71.880 ;
        RECT 23.470 66.460 23.850 69.480 ;
        RECT 25.650 68.910 25.930 71.315 ;
        RECT 26.260 67.755 26.560 74.795 ;
        RECT 27.380 67.150 27.680 74.080 ;
        RECT 28.690 67.750 28.990 74.100 ;
        RECT 29.285 69.625 29.610 74.785 ;
        RECT 30.005 67.780 30.300 74.605 ;
        RECT 31.135 67.240 31.435 74.050 ;
        RECT 31.925 67.835 32.235 74.025 ;
        RECT 32.720 67.765 33.020 74.595 ;
        RECT 33.845 67.150 34.145 74.090 ;
        RECT 35.295 67.025 35.575 70.060 ;
        RECT 36.055 67.725 36.375 74.085 ;
        RECT 36.905 67.725 37.205 74.545 ;
        RECT 38.045 66.980 38.345 74.135 ;
        RECT 38.680 69.125 39.060 69.505 ;
        RECT 39.385 65.010 39.745 71.570 ;
        RECT 40.525 69.760 40.850 71.625 ;
        RECT 41.190 66.415 41.650 71.100 ;
        RECT 41.975 68.960 42.425 77.780 ;
        RECT 44.160 70.785 44.590 73.775 ;
        RECT 41.905 65.070 42.285 65.450 ;
        RECT 44.795 65.090 45.175 66.465 ;
        RECT 45.565 65.910 45.880 76.960 ;
        RECT 46.580 75.655 46.870 77.715 ;
        RECT 46.500 67.800 46.825 70.170 ;
        RECT 48.150 69.845 48.550 73.810 ;
        RECT 48.870 65.740 49.195 68.505 ;
        RECT 49.855 67.775 50.260 71.105 ;
        RECT 54.505 64.800 54.875 73.900 ;
        RECT 55.450 65.865 55.740 77.700 ;
        RECT 63.355 75.595 63.665 78.110 ;
        RECT 59.265 67.830 59.705 71.105 ;
        RECT 61.645 69.845 62.170 73.785 ;
        RECT 60.805 65.740 61.130 68.505 ;
        RECT 63.320 67.835 63.735 70.225 ;
        RECT 64.350 66.395 64.665 77.080 ;
        RECT 65.680 70.785 66.165 73.795 ;
        RECT 65.050 65.005 65.385 66.355 ;
        RECT 4.770 49.035 5.125 62.945 ;
        RECT 68.115 62.315 68.565 72.580 ;
        RECT 6.395 49.955 6.755 61.345 ;
        RECT 69.280 60.775 69.765 69.660 ;
        RECT 76.110 60.130 76.515 72.010 ;
        RECT 78.185 62.030 78.575 73.610 ;
        RECT 81.455 65.950 81.810 77.035 ;
        RECT 85.200 75.675 85.490 77.735 ;
        RECT 91.980 74.525 92.290 74.555 ;
        RECT 82.780 70.805 83.250 73.795 ;
        RECT 85.130 67.820 85.445 70.190 ;
        RECT 86.750 69.865 87.170 73.830 ;
        RECT 83.415 65.110 83.795 66.485 ;
        RECT 87.490 65.760 87.815 68.525 ;
        RECT 88.475 67.795 88.880 71.125 ;
        RECT 91.980 68.425 92.295 74.525 ;
        RECT 93.125 64.820 93.495 73.920 ;
        RECT 94.070 65.885 94.360 77.720 ;
        RECT 101.975 75.615 102.285 78.130 ;
        RECT 106.225 77.315 106.605 77.695 ;
        RECT 108.355 77.315 108.735 77.695 ;
        RECT 94.965 68.380 95.295 74.575 ;
        RECT 97.870 67.850 98.325 71.125 ;
        RECT 100.230 69.865 100.775 73.805 ;
        RECT 104.285 70.805 104.720 73.815 ;
        RECT 99.425 65.760 99.750 68.525 ;
        RECT 101.940 67.855 102.355 70.245 ;
        RECT 105.480 66.430 105.810 77.125 ;
        RECT 106.915 70.765 107.300 76.550 ;
        RECT 103.670 65.025 104.005 66.375 ;
        RECT 107.275 66.010 107.700 70.285 ;
        RECT 108.975 67.775 109.275 74.815 ;
        RECT 110.095 67.170 110.395 74.100 ;
        RECT 111.405 67.770 111.705 74.120 ;
        RECT 105.935 65.100 106.315 65.480 ;
        RECT 108.130 65.085 108.510 65.465 ;
        RECT 112.000 65.025 112.290 74.805 ;
        RECT 112.720 67.800 113.015 74.625 ;
        RECT 113.850 67.260 114.150 74.070 ;
        RECT 114.640 67.855 114.950 77.895 ;
        RECT 123.830 76.140 124.210 76.520 ;
        RECT 115.435 67.785 115.735 74.615 ;
        RECT 116.560 67.170 116.860 74.110 ;
        RECT 118.010 67.045 118.290 70.080 ;
        RECT 118.770 67.745 119.050 74.105 ;
        RECT 119.620 67.745 119.920 74.565 ;
        RECT 120.760 67.000 121.060 74.155 ;
        RECT 121.405 71.190 121.785 71.570 ;
        RECT 121.405 69.135 121.785 69.515 ;
        RECT 123.255 69.015 123.570 73.340 ;
        RECT 123.865 71.090 124.145 72.620 ;
        RECT 124.435 67.775 124.735 74.815 ;
        RECT 126.210 68.530 126.510 72.590 ;
        RECT 123.730 65.965 124.110 66.345 ;
        RECT 127.460 65.560 127.750 74.805 ;
        RECT 129.310 67.260 129.610 74.070 ;
        RECT 130.100 67.855 130.410 76.590 ;
        RECT 130.895 67.785 131.195 74.615 ;
        RECT 132.700 68.515 132.980 72.605 ;
        RECT 133.470 67.045 133.750 70.080 ;
        RECT 136.220 67.000 136.520 74.155 ;
        RECT 138.300 72.875 138.675 81.155 ;
        RECT 140.045 72.035 140.345 83.145 ;
        RECT 11.870 47.340 12.170 54.270 ;
        RECT 13.180 47.940 13.480 54.290 ;
        RECT 14.495 47.970 14.790 54.795 ;
        RECT 18.335 47.340 18.635 54.280 ;
        RECT 20.545 47.915 20.850 54.275 ;
        RECT 21.395 47.915 21.695 54.735 ;
        RECT 23.205 51.360 23.585 51.740 ;
        RECT 24.990 49.940 25.310 52.070 ;
        RECT 23.420 46.650 23.800 49.670 ;
        RECT 25.600 49.100 25.880 51.505 ;
        RECT 26.210 47.945 26.510 54.985 ;
        RECT 27.330 47.340 27.630 54.270 ;
        RECT 28.640 47.940 28.940 54.290 ;
        RECT 29.235 49.815 29.560 54.975 ;
        RECT 29.955 47.970 30.250 54.795 ;
        RECT 31.085 47.430 31.385 54.240 ;
        RECT 31.875 48.025 32.185 54.215 ;
        RECT 32.670 47.955 32.970 54.785 ;
        RECT 33.795 47.340 34.095 54.280 ;
        RECT 35.245 47.215 35.525 50.250 ;
        RECT 36.005 47.915 36.325 54.275 ;
        RECT 36.855 47.915 37.155 54.735 ;
        RECT 37.995 47.170 38.295 54.325 ;
        RECT 38.630 49.315 39.010 49.695 ;
        RECT 39.335 45.200 39.695 51.760 ;
        RECT 40.475 49.950 40.800 51.815 ;
        RECT 41.140 46.605 41.600 51.290 ;
        RECT 41.925 49.150 42.375 57.970 ;
        RECT 44.110 50.975 44.540 53.965 ;
        RECT 41.855 45.260 42.235 45.640 ;
        RECT 44.745 45.280 45.125 46.655 ;
        RECT 45.515 46.100 45.830 57.150 ;
        RECT 46.530 55.845 46.820 57.905 ;
        RECT 46.450 47.990 46.775 50.360 ;
        RECT 48.100 50.035 48.500 54.000 ;
        RECT 48.820 45.930 49.145 48.695 ;
        RECT 49.805 47.965 50.210 51.295 ;
        RECT 54.455 44.990 54.825 54.090 ;
        RECT 55.400 46.055 55.690 57.890 ;
        RECT 63.305 55.785 63.615 58.300 ;
        RECT 59.215 48.020 59.655 51.295 ;
        RECT 61.595 50.035 62.120 53.975 ;
        RECT 60.755 45.930 61.080 48.695 ;
        RECT 63.270 48.025 63.685 50.415 ;
        RECT 64.300 46.585 64.615 57.270 ;
        RECT 65.630 50.975 66.115 53.985 ;
        RECT 65.000 45.195 65.335 46.545 ;
        RECT 4.770 29.195 5.125 43.135 ;
        RECT 68.115 42.505 68.565 52.770 ;
        RECT 6.395 29.985 6.755 41.535 ;
        RECT 69.280 40.965 69.765 49.850 ;
        RECT 76.220 40.240 76.625 52.285 ;
        RECT 78.295 42.140 78.685 53.565 ;
        RECT 81.455 45.980 81.810 57.065 ;
        RECT 85.200 55.705 85.490 57.765 ;
        RECT 91.980 54.555 92.290 54.585 ;
        RECT 82.780 50.835 83.250 53.825 ;
        RECT 85.130 47.850 85.445 50.220 ;
        RECT 86.750 49.895 87.170 53.860 ;
        RECT 83.415 45.140 83.795 46.515 ;
        RECT 87.490 45.790 87.815 48.555 ;
        RECT 88.475 47.825 88.880 51.155 ;
        RECT 91.980 48.455 92.295 54.555 ;
        RECT 93.125 44.850 93.495 53.950 ;
        RECT 94.070 45.915 94.360 57.750 ;
        RECT 101.975 55.645 102.285 58.160 ;
        RECT 106.225 57.345 106.605 57.725 ;
        RECT 108.355 57.345 108.735 57.725 ;
        RECT 94.965 48.410 95.295 54.605 ;
        RECT 97.870 47.880 98.325 51.155 ;
        RECT 100.230 49.895 100.775 53.835 ;
        RECT 104.285 50.835 104.720 53.845 ;
        RECT 99.425 45.790 99.750 48.555 ;
        RECT 101.940 47.885 102.355 50.275 ;
        RECT 105.480 46.460 105.810 57.155 ;
        RECT 106.915 50.795 107.300 56.580 ;
        RECT 103.670 45.055 104.005 46.405 ;
        RECT 107.275 46.040 107.700 50.315 ;
        RECT 108.975 47.805 109.275 54.845 ;
        RECT 110.095 47.200 110.395 54.130 ;
        RECT 111.405 47.800 111.705 54.150 ;
        RECT 105.935 45.130 106.315 45.510 ;
        RECT 108.130 45.115 108.510 45.495 ;
        RECT 112.000 45.055 112.290 54.835 ;
        RECT 112.720 47.830 113.015 54.655 ;
        RECT 113.850 47.290 114.150 54.100 ;
        RECT 114.640 47.885 114.950 57.925 ;
        RECT 123.830 56.170 124.210 56.550 ;
        RECT 115.435 47.815 115.735 54.645 ;
        RECT 116.560 47.200 116.860 54.140 ;
        RECT 118.010 47.075 118.290 50.110 ;
        RECT 118.770 47.775 119.050 54.135 ;
        RECT 119.620 47.775 119.920 54.595 ;
        RECT 120.760 47.030 121.060 54.185 ;
        RECT 121.405 51.220 121.785 51.600 ;
        RECT 121.405 49.165 121.785 49.545 ;
        RECT 123.255 49.045 123.570 53.370 ;
        RECT 123.865 51.120 124.145 52.650 ;
        RECT 124.435 47.805 124.735 54.845 ;
        RECT 126.210 48.560 126.510 52.620 ;
        RECT 123.730 45.995 124.110 46.375 ;
        RECT 127.460 45.590 127.750 54.835 ;
        RECT 129.310 47.290 129.610 54.100 ;
        RECT 130.100 47.885 130.410 56.620 ;
        RECT 130.895 47.815 131.195 54.645 ;
        RECT 132.700 48.545 132.980 52.635 ;
        RECT 133.470 47.075 133.750 50.110 ;
        RECT 136.220 47.030 136.520 54.185 ;
        RECT 138.560 52.800 138.935 61.000 ;
        RECT 140.305 51.995 140.605 62.990 ;
        RECT 11.840 27.545 12.140 34.475 ;
        RECT 13.150 28.145 13.450 34.495 ;
        RECT 14.465 28.175 14.760 35.000 ;
        RECT 18.305 27.545 18.605 34.485 ;
        RECT 20.515 28.120 20.820 34.480 ;
        RECT 21.365 28.120 21.665 34.940 ;
        RECT 23.175 31.565 23.555 31.945 ;
        RECT 24.960 30.145 25.280 32.275 ;
        RECT 23.390 26.855 23.770 29.875 ;
        RECT 25.570 29.305 25.850 31.710 ;
        RECT 26.180 28.150 26.480 35.190 ;
        RECT 27.300 27.545 27.600 34.475 ;
        RECT 28.610 28.145 28.910 34.495 ;
        RECT 29.205 30.020 29.530 35.180 ;
        RECT 29.925 28.175 30.220 35.000 ;
        RECT 31.055 27.635 31.355 34.445 ;
        RECT 31.845 28.230 32.155 34.420 ;
        RECT 32.640 28.160 32.940 34.990 ;
        RECT 33.765 27.545 34.065 34.485 ;
        RECT 35.215 27.420 35.495 30.455 ;
        RECT 35.975 28.120 36.295 34.480 ;
        RECT 36.825 28.120 37.125 34.940 ;
        RECT 37.965 27.375 38.265 34.530 ;
        RECT 38.600 29.520 38.980 29.900 ;
        RECT 39.305 25.405 39.665 31.965 ;
        RECT 40.445 30.155 40.770 32.020 ;
        RECT 41.110 26.810 41.570 31.495 ;
        RECT 41.895 29.355 42.345 38.175 ;
        RECT 44.080 31.180 44.510 34.170 ;
        RECT 41.825 25.465 42.205 25.845 ;
        RECT 44.715 25.485 45.095 26.860 ;
        RECT 45.485 26.305 45.800 37.355 ;
        RECT 46.500 36.050 46.790 38.110 ;
        RECT 46.420 28.195 46.745 30.565 ;
        RECT 48.070 30.240 48.470 34.205 ;
        RECT 48.790 26.135 49.115 28.900 ;
        RECT 49.775 28.170 50.180 31.500 ;
        RECT 54.425 25.195 54.795 34.295 ;
        RECT 55.370 26.260 55.660 38.095 ;
        RECT 63.275 35.990 63.585 38.505 ;
        RECT 59.185 28.225 59.625 31.500 ;
        RECT 61.565 30.240 62.090 34.180 ;
        RECT 60.725 26.135 61.050 28.900 ;
        RECT 63.240 28.230 63.655 30.620 ;
        RECT 64.270 26.790 64.585 37.475 ;
        RECT 65.600 31.180 66.085 34.190 ;
        RECT 72.060 33.100 75.385 33.690 ;
        RECT 72.060 32.485 72.810 33.100 ;
        RECT 73.965 29.645 74.635 32.295 ;
        RECT 64.970 25.400 65.305 26.750 ;
        RECT 75.925 13.490 76.375 32.530 ;
        RECT 77.715 12.715 78.130 33.895 ;
        RECT 81.455 26.315 81.810 37.400 ;
        RECT 85.200 36.040 85.490 38.100 ;
        RECT 91.980 34.890 92.290 34.920 ;
        RECT 82.780 31.170 83.250 34.160 ;
        RECT 85.130 28.185 85.445 30.555 ;
        RECT 86.750 30.230 87.170 34.195 ;
        RECT 83.415 25.475 83.795 26.850 ;
        RECT 87.490 26.125 87.815 28.890 ;
        RECT 88.475 28.160 88.880 31.490 ;
        RECT 91.980 28.790 92.295 34.890 ;
        RECT 93.125 25.185 93.495 34.285 ;
        RECT 94.070 26.250 94.360 38.085 ;
        RECT 101.975 35.980 102.285 38.495 ;
        RECT 106.225 37.680 106.605 38.060 ;
        RECT 108.355 37.680 108.735 38.060 ;
        RECT 94.965 28.745 95.295 34.940 ;
        RECT 97.870 28.215 98.325 31.490 ;
        RECT 100.230 30.230 100.775 34.170 ;
        RECT 104.285 31.170 104.720 34.180 ;
        RECT 99.425 26.125 99.750 28.890 ;
        RECT 101.940 28.220 102.355 30.610 ;
        RECT 105.480 26.795 105.810 37.490 ;
        RECT 106.915 31.130 107.300 36.915 ;
        RECT 103.670 25.390 104.005 26.740 ;
        RECT 107.275 26.375 107.700 30.650 ;
        RECT 108.975 28.140 109.275 35.180 ;
        RECT 110.095 27.535 110.395 34.465 ;
        RECT 111.405 28.135 111.705 34.485 ;
        RECT 105.935 25.465 106.315 25.845 ;
        RECT 108.130 25.450 108.510 25.830 ;
        RECT 112.000 25.390 112.290 35.170 ;
        RECT 112.720 28.165 113.015 34.990 ;
        RECT 113.850 27.625 114.150 34.435 ;
        RECT 114.640 28.220 114.950 38.260 ;
        RECT 123.830 36.505 124.210 36.885 ;
        RECT 115.435 28.150 115.735 34.980 ;
        RECT 116.560 27.535 116.860 34.475 ;
        RECT 118.010 27.410 118.290 30.445 ;
        RECT 118.770 28.110 119.050 34.470 ;
        RECT 119.620 28.110 119.920 34.930 ;
        RECT 120.760 27.365 121.060 34.520 ;
        RECT 121.405 31.555 121.785 31.935 ;
        RECT 121.405 29.500 121.785 29.880 ;
        RECT 123.255 29.380 123.570 33.705 ;
        RECT 123.865 31.455 124.145 32.985 ;
        RECT 124.435 28.140 124.735 35.180 ;
        RECT 126.210 28.895 126.510 32.955 ;
        RECT 123.730 26.330 124.110 26.710 ;
        RECT 127.460 25.925 127.750 35.170 ;
        RECT 129.310 27.625 129.610 34.435 ;
        RECT 130.100 28.220 130.410 36.955 ;
        RECT 130.895 28.150 131.195 34.980 ;
        RECT 132.700 28.880 132.980 32.970 ;
        RECT 133.470 27.410 133.750 30.445 ;
        RECT 136.220 27.365 136.520 34.520 ;
        RECT 138.145 33.285 138.520 41.125 ;
        RECT 140.000 32.535 140.300 43.075 ;
        RECT 82.130 9.160 82.430 13.220 ;
        RECT 88.620 9.145 88.900 13.235 ;
      LAYER Metal3 ;
        RECT 106.180 334.030 108.775 334.460 ;
        RECT 106.860 332.905 124.230 333.245 ;
        RECT 23.235 328.015 40.960 328.335 ;
        RECT 38.650 325.895 42.550 326.380 ;
        RECT 23.400 323.240 41.700 323.625 ;
        RECT 107.115 322.705 124.300 323.190 ;
        RECT 39.280 321.920 42.345 322.245 ;
        RECT 105.925 321.790 108.520 322.240 ;
        RECT 4.710 319.165 68.590 319.585 ;
        RECT 77.265 319.290 140.710 319.910 ;
        RECT 6.350 317.620 69.790 318.110 ;
        RECT 75.170 317.335 138.895 317.905 ;
        RECT 105.980 314.305 108.575 314.735 ;
        RECT 106.660 313.180 124.030 313.520 ;
        RECT 23.190 308.325 40.915 308.645 ;
        RECT 121.185 308.210 124.030 308.590 ;
        RECT 4.705 306.950 25.410 307.245 ;
        RECT 4.525 306.085 25.995 306.380 ;
        RECT 38.605 306.205 42.505 306.690 ;
        RECT 121.160 306.135 123.445 306.560 ;
        RECT 23.355 303.550 41.655 303.935 ;
        RECT 106.915 302.980 124.100 303.465 ;
        RECT 39.235 302.230 42.300 302.555 ;
        RECT 105.725 302.065 108.320 302.515 ;
        RECT 4.710 299.665 68.590 300.085 ;
        RECT 77.565 299.540 141.010 300.160 ;
        RECT 6.350 298.120 69.790 298.610 ;
        RECT 75.470 297.585 139.195 298.155 ;
        RECT 106.135 294.660 108.730 295.090 ;
        RECT 106.815 293.535 124.185 293.875 ;
        RECT 23.380 288.615 41.105 288.935 ;
        RECT 121.340 288.565 124.185 288.945 ;
        RECT 4.895 287.240 25.600 287.535 ;
        RECT 4.715 286.375 26.185 286.670 ;
        RECT 38.795 286.495 42.695 286.980 ;
        RECT 121.315 286.490 123.600 286.915 ;
        RECT 23.545 283.840 41.845 284.225 ;
        RECT 107.070 283.335 124.255 283.820 ;
        RECT 39.425 282.520 42.490 282.845 ;
        RECT 105.880 282.420 108.475 282.870 ;
        RECT 4.920 279.625 68.800 280.045 ;
        RECT 77.585 279.880 141.030 280.500 ;
        RECT 6.560 278.080 70.000 278.570 ;
        RECT 75.490 277.925 139.215 278.495 ;
        RECT 106.135 274.865 108.730 275.295 ;
        RECT 106.815 273.740 124.185 274.080 ;
        RECT 23.185 268.775 40.910 269.095 ;
        RECT 121.340 268.770 124.185 269.150 ;
        RECT 4.700 267.400 25.405 267.695 ;
        RECT 4.520 266.535 25.990 266.830 ;
        RECT 38.600 266.655 42.500 267.140 ;
        RECT 121.315 266.695 123.600 267.120 ;
        RECT 23.350 264.000 41.650 264.385 ;
        RECT 107.070 263.540 124.255 264.025 ;
        RECT 39.230 262.680 42.295 263.005 ;
        RECT 105.880 262.625 108.475 263.075 ;
        RECT 4.875 259.835 68.755 260.255 ;
        RECT 77.585 260.145 141.030 260.765 ;
        RECT 6.515 258.290 69.955 258.780 ;
        RECT 75.490 258.190 139.215 258.760 ;
        RECT 106.055 255.110 108.650 255.540 ;
        RECT 106.735 253.985 124.105 254.325 ;
        RECT 23.055 249.065 40.780 249.385 ;
        RECT 121.260 249.015 124.105 249.395 ;
        RECT 4.570 247.690 25.275 247.985 ;
        RECT 4.390 246.825 25.860 247.120 ;
        RECT 38.470 246.945 42.370 247.430 ;
        RECT 121.235 246.940 123.520 247.365 ;
        RECT 23.220 244.290 41.520 244.675 ;
        RECT 106.990 243.785 124.175 244.270 ;
        RECT 39.100 242.970 42.165 243.295 ;
        RECT 105.800 242.870 108.395 243.320 ;
        RECT 4.570 240.205 68.450 240.625 ;
        RECT 77.485 240.440 140.930 241.060 ;
        RECT 6.210 238.660 69.650 239.150 ;
        RECT 75.390 238.485 139.115 239.055 ;
        RECT 106.160 235.395 108.755 235.825 ;
        RECT 106.840 234.270 124.210 234.610 ;
        RECT 23.185 229.305 40.910 229.625 ;
        RECT 121.365 229.300 124.210 229.680 ;
        RECT 4.700 227.930 25.405 228.225 ;
        RECT 4.520 227.065 25.990 227.360 ;
        RECT 38.600 227.185 42.500 227.670 ;
        RECT 121.340 227.225 123.625 227.650 ;
        RECT 23.350 224.530 41.650 224.915 ;
        RECT 107.095 224.070 124.280 224.555 ;
        RECT 39.230 223.210 42.295 223.535 ;
        RECT 105.905 223.155 108.500 223.605 ;
        RECT 4.665 220.430 68.545 220.850 ;
        RECT 77.745 220.285 141.190 220.905 ;
        RECT 6.305 218.885 69.745 219.375 ;
        RECT 75.650 218.330 139.375 218.900 ;
        RECT 106.160 215.425 108.755 215.855 ;
        RECT 106.840 214.300 124.210 214.640 ;
        RECT 23.135 209.495 40.860 209.815 ;
        RECT 121.365 209.330 124.210 209.710 ;
        RECT 4.650 208.120 25.355 208.415 ;
        RECT 4.470 207.255 25.940 207.550 ;
        RECT 38.550 207.375 42.450 207.860 ;
        RECT 121.340 207.255 123.625 207.680 ;
        RECT 23.300 204.720 41.600 205.105 ;
        RECT 107.095 204.100 124.280 204.585 ;
        RECT 39.180 203.400 42.245 203.725 ;
        RECT 105.905 203.185 108.500 203.635 ;
        RECT 4.665 200.620 68.545 201.040 ;
        RECT 77.855 200.395 141.300 201.015 ;
        RECT 6.305 199.075 69.745 199.565 ;
        RECT 75.760 198.440 139.485 199.010 ;
        RECT 106.160 195.760 108.755 196.190 ;
        RECT 106.840 194.635 124.210 194.975 ;
        RECT 23.105 189.700 40.830 190.020 ;
        RECT 121.365 189.665 124.210 190.045 ;
        RECT 4.620 188.325 25.325 188.620 ;
        RECT 4.440 187.460 25.910 187.755 ;
        RECT 38.520 187.580 42.420 188.065 ;
        RECT 121.340 187.590 123.625 188.015 ;
        RECT 23.270 184.925 41.570 185.310 ;
        RECT 107.095 184.435 124.280 184.920 ;
        RECT 39.150 183.605 42.215 183.930 ;
        RECT 105.905 183.520 108.500 183.970 ;
        RECT 4.505 180.435 69.155 180.920 ;
        RECT 77.225 180.705 141.010 181.335 ;
        RECT 6.450 179.060 70.860 179.600 ;
        RECT 75.295 179.410 139.280 179.945 ;
        RECT 106.200 175.920 108.795 176.350 ;
        RECT 106.880 174.795 124.250 175.135 ;
        RECT 23.255 169.905 40.980 170.225 ;
        RECT 121.405 169.825 124.250 170.205 ;
        RECT 4.770 168.530 25.475 168.825 ;
        RECT 4.590 167.665 26.060 167.960 ;
        RECT 38.670 167.785 42.570 168.270 ;
        RECT 121.380 167.750 123.665 168.175 ;
        RECT 23.420 165.130 41.720 165.515 ;
        RECT 107.135 164.595 124.320 165.080 ;
        RECT 39.300 163.810 42.365 164.135 ;
        RECT 105.945 163.680 108.540 164.130 ;
        RECT 4.730 161.055 68.610 161.475 ;
        RECT 77.285 161.180 140.730 161.800 ;
        RECT 6.370 159.510 69.810 160.000 ;
        RECT 75.190 159.225 138.915 159.795 ;
        RECT 106.000 156.195 108.595 156.625 ;
        RECT 106.680 155.070 124.050 155.410 ;
        RECT 23.210 150.215 40.935 150.535 ;
        RECT 121.205 150.100 124.050 150.480 ;
        RECT 4.725 148.840 25.430 149.135 ;
        RECT 4.545 147.975 26.015 148.270 ;
        RECT 38.625 148.095 42.525 148.580 ;
        RECT 121.180 148.025 123.465 148.450 ;
        RECT 23.375 145.440 41.675 145.825 ;
        RECT 106.935 144.870 124.120 145.355 ;
        RECT 39.255 144.120 42.320 144.445 ;
        RECT 105.745 143.955 108.340 144.405 ;
        RECT 4.730 141.555 68.610 141.975 ;
        RECT 77.585 141.430 141.030 142.050 ;
        RECT 6.370 140.010 69.810 140.500 ;
        RECT 75.490 139.475 139.215 140.045 ;
        RECT 106.155 136.550 108.750 136.980 ;
        RECT 106.835 135.425 124.205 135.765 ;
        RECT 23.400 130.505 41.125 130.825 ;
        RECT 121.360 130.455 124.205 130.835 ;
        RECT 4.915 129.130 25.620 129.425 ;
        RECT 4.735 128.265 26.205 128.560 ;
        RECT 38.815 128.385 42.715 128.870 ;
        RECT 121.335 128.380 123.620 128.805 ;
        RECT 23.565 125.730 41.865 126.115 ;
        RECT 107.090 125.225 124.275 125.710 ;
        RECT 39.445 124.410 42.510 124.735 ;
        RECT 105.900 124.310 108.495 124.760 ;
        RECT 4.940 121.515 68.820 121.935 ;
        RECT 77.605 121.770 141.050 122.390 ;
        RECT 6.580 119.970 70.020 120.460 ;
        RECT 75.510 119.815 139.235 120.385 ;
        RECT 106.155 116.755 108.750 117.185 ;
        RECT 106.835 115.630 124.205 115.970 ;
        RECT 23.205 110.665 40.930 110.985 ;
        RECT 121.360 110.660 124.205 111.040 ;
        RECT 4.720 109.290 25.425 109.585 ;
        RECT 4.540 108.425 26.010 108.720 ;
        RECT 38.620 108.545 42.520 109.030 ;
        RECT 121.335 108.585 123.620 109.010 ;
        RECT 23.370 105.890 41.670 106.275 ;
        RECT 107.090 105.430 124.275 105.915 ;
        RECT 39.250 104.570 42.315 104.895 ;
        RECT 105.900 104.515 108.495 104.965 ;
        RECT 4.895 101.725 68.775 102.145 ;
        RECT 77.605 102.035 141.050 102.655 ;
        RECT 6.535 100.180 69.975 100.670 ;
        RECT 75.510 100.080 139.235 100.650 ;
        RECT 106.075 97.000 108.670 97.430 ;
        RECT 106.755 95.875 124.125 96.215 ;
        RECT 23.075 90.955 40.800 91.275 ;
        RECT 121.280 90.905 124.125 91.285 ;
        RECT 4.590 89.580 25.295 89.875 ;
        RECT 4.410 88.715 25.880 89.010 ;
        RECT 38.490 88.835 42.390 89.320 ;
        RECT 121.255 88.830 123.540 89.255 ;
        RECT 23.240 86.180 41.540 86.565 ;
        RECT 107.010 85.675 124.195 86.160 ;
        RECT 39.120 84.860 42.185 85.185 ;
        RECT 105.820 84.760 108.415 85.210 ;
        RECT 4.590 82.095 68.470 82.515 ;
        RECT 77.505 82.330 140.950 82.950 ;
        RECT 6.230 80.550 69.670 81.040 ;
        RECT 75.410 80.375 139.135 80.945 ;
        RECT 106.180 77.285 108.775 77.715 ;
        RECT 106.860 76.160 124.230 76.500 ;
        RECT 23.205 71.195 40.930 71.515 ;
        RECT 121.385 71.190 124.230 71.570 ;
        RECT 4.720 69.820 25.425 70.115 ;
        RECT 4.540 68.955 26.010 69.250 ;
        RECT 38.620 69.075 42.520 69.560 ;
        RECT 121.360 69.115 123.645 69.540 ;
        RECT 23.370 66.420 41.670 66.805 ;
        RECT 107.115 65.960 124.300 66.445 ;
        RECT 39.250 65.100 42.315 65.425 ;
        RECT 105.925 65.045 108.520 65.495 ;
        RECT 4.685 62.320 68.565 62.740 ;
        RECT 77.765 62.175 141.210 62.795 ;
        RECT 6.325 60.775 69.765 61.265 ;
        RECT 75.670 60.220 139.395 60.790 ;
        RECT 106.180 57.315 108.775 57.745 ;
        RECT 106.860 56.190 124.230 56.530 ;
        RECT 23.155 51.385 40.880 51.705 ;
        RECT 121.385 51.220 124.230 51.600 ;
        RECT 4.670 50.010 25.375 50.305 ;
        RECT 4.490 49.145 25.960 49.440 ;
        RECT 38.570 49.265 42.470 49.750 ;
        RECT 121.360 49.145 123.645 49.570 ;
        RECT 23.320 46.610 41.620 46.995 ;
        RECT 107.115 45.990 124.300 46.475 ;
        RECT 39.200 45.290 42.265 45.615 ;
        RECT 105.925 45.075 108.520 45.525 ;
        RECT 4.685 42.510 68.565 42.930 ;
        RECT 77.875 42.285 141.320 42.905 ;
        RECT 6.325 40.965 69.765 41.455 ;
        RECT 75.780 40.330 139.505 40.900 ;
        RECT 106.180 37.650 108.775 38.080 ;
        RECT 106.860 36.525 124.230 36.865 ;
        RECT 23.125 31.590 40.850 31.910 ;
        RECT 121.385 31.555 124.230 31.935 ;
        RECT 4.640 30.215 25.345 30.510 ;
        RECT 4.460 29.350 25.930 29.645 ;
        RECT 38.540 29.470 42.440 29.955 ;
        RECT 121.360 29.480 123.645 29.905 ;
        RECT 23.290 26.815 41.590 27.200 ;
        RECT 107.115 26.325 124.300 26.810 ;
        RECT 39.170 25.495 42.235 25.820 ;
        RECT 105.925 25.410 108.520 25.860 ;
  END
END fa16b_rev
END LIBRARY

