`default_nettype none

(* blackbox *)
module fa8b_rev (
    inout wire z,
    inout wire z_not,
    inout wire c0_b,
    inout wire c0_not_b,
    inout wire c7_not,
    inout wire c7,
    inout wire s5_not,
    inout wire s5,
    inout wire s0_not,
    inout wire s0,
    inout wire s6_not,
    inout wire s6,
    inout wire s1_not,
    inout wire s1,
    inout wire s7_not,
    inout wire s7,
    inout wire s2_not,
    inout wire s2,
    inout wire s3_not,
    inout wire s3,
    inout wire s4_not,
    inout wire s4,
    inout wire c0_f,
    inout wire c0_f_not,
    inout wire VSS,
    inout wire VDD,
    inout wire a0_f,
    inout wire a0_not_f,
    inout wire b0,
    inout wire b0_not,
    inout wire a1_f,
    inout wire a1_not_f,
    inout wire b1,
    inout wire b1_not,
    inout wire a2_f,
    inout wire a2_not_f,
    inout wire b2,
    inout wire b2_not,
    inout wire a3_f,
    inout wire a3_not_f,
    inout wire b3,
    inout wire b3_not,
    inout wire a4_f,
    inout wire a4_not_f,
    inout wire b4,
    inout wire b4_not,
    inout wire a5_f,
    inout wire a5_not_f,
    inout wire b5,
    inout wire b5_not,
    inout wire a6_f,
    inout wire a6_not_f,
    inout wire b6,
    inout wire b6_not,
    inout wire a7_f,
    inout wire a7_not_f,
    inout wire b7,
    inout wire b7_not,
    inout wire a0_b,
    inout wire a0_not_b,
    inout wire a1_b,
    inout wire a1_not_b,
    inout wire a2_b,
    inout wire a2_not_b,
    inout wire a3_b,
    inout wire a3_not_b,
    inout wire a4_b,
    inout wire a4_not_b,
    inout wire a5_b,
    inout wire a5_not_b,
    inout wire a6_b,
    inout wire a6_not_b,
    inout wire a7_b,
    inout wire a7_not_b
);

endmodule
