VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO 16b_FA
  CLASS BLOCK ;
  FOREIGN 16b_FA ;
  ORIGIN 0.000 0.000 ;
  SIZE 169.925 BY 349.940 ;
  PIN vss
    ANTENNADIFFAREA 36.745197 ;
    PORT
      LAYER Metal3 ;
        RECT 153.995 322.695 156.130 323.595 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 153.995 302.925 156.130 303.825 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 153.995 283.230 156.130 284.130 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 153.995 263.495 156.130 264.395 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 153.995 243.740 156.130 244.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 154.015 223.990 156.150 224.890 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 154.015 204.045 156.150 204.945 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 153.995 184.350 156.130 185.250 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 10.275 243.740 81.245 244.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 10.275 283.230 81.245 284.130 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 10.295 223.990 81.265 224.890 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 10.275 302.925 81.245 303.825 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 10.295 204.045 81.265 204.945 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 10.275 263.495 81.245 264.395 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 10.275 184.350 81.245 185.250 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 10.275 322.695 81.245 323.595 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 10.330 164.580 81.300 165.480 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 10.275 144.845 81.245 145.745 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 10.275 125.165 81.245 126.065 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 10.295 105.375 81.265 106.275 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 10.310 85.595 81.280 86.495 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 10.215 65.865 81.185 66.765 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 10.310 45.910 81.280 46.810 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 10.325 26.285 81.295 27.185 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 10.290 6.510 81.260 7.410 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 153.995 144.845 156.130 145.745 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 154.030 45.910 156.165 46.810 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 154.015 105.375 156.150 106.275 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 154.045 26.285 156.180 27.185 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 154.050 164.580 156.185 165.480 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 154.010 6.510 156.145 7.410 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 154.030 85.595 156.165 86.495 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 153.995 125.165 156.130 126.065 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 153.935 65.865 156.070 66.765 ;
    END
  END vss
  PIN vdd
    ANTENNADIFFAREA 59.785198 ;
    PORT
      LAYER Metal3 ;
        RECT 155.735 179.540 156.140 180.440 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 155.735 199.380 156.140 200.280 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 155.755 219.065 156.160 219.965 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 155.720 239.030 156.125 239.930 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 155.755 258.740 156.160 259.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 155.745 278.490 156.150 279.390 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 155.735 298.285 156.140 299.185 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 155.745 317.925 156.150 318.825 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 155.740 337.670 156.145 338.570 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9.630 199.380 11.810 200.280 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9.650 219.065 11.830 219.965 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9.615 239.030 11.795 239.930 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9.650 258.740 11.830 259.640 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9.640 278.490 11.820 279.390 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9.630 298.285 11.810 299.185 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9.640 317.925 11.820 318.825 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9.635 337.670 11.815 338.570 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9.630 179.540 11.810 180.440 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9.630 21.560 11.810 22.460 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9.645 41.340 11.825 42.240 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9.665 60.980 11.845 61.880 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9.630 80.910 11.810 81.810 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9.630 100.650 11.810 101.550 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9.630 120.340 11.810 121.240 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9.640 140.180 11.820 141.080 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9.640 159.845 11.820 160.745 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 155.770 60.980 156.175 61.880 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 155.735 80.910 156.140 81.810 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 155.735 100.650 156.140 101.550 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 155.735 120.340 156.140 121.240 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 155.745 140.180 156.150 141.080 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 155.745 159.845 156.150 160.745 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 155.735 21.560 156.140 22.460 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 155.750 41.340 156.155 42.240 ;
    END
  END vdd
  PIN c0_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal3 ;
        RECT 149.280 332.675 151.215 332.985 ;
    END
  END c0_b
  PIN a0_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 132.195 336.890 147.930 337.300 ;
    END
  END a0_b
  PIN a0_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 132.790 336.110 147.920 336.565 ;
    END
  END a0_not_b
  PIN a1_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 131.995 317.165 147.730 317.575 ;
    END
  END a1_b
  PIN a1_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 132.590 316.385 147.720 316.840 ;
    END
  END a1_not_b
  PIN a2_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 132.150 297.520 147.885 297.930 ;
    END
  END a2_b
  PIN a2_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 132.745 296.740 147.875 297.195 ;
    END
  END a2_not_b
  PIN a3_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 132.150 277.725 147.885 278.135 ;
    END
  END a3_b
  PIN a3_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 132.745 276.945 147.875 277.400 ;
    END
  END a3_not_b
  PIN a4_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 132.070 257.970 147.805 258.380 ;
    END
  END a4_b
  PIN a4_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 132.665 257.190 147.795 257.645 ;
    END
  END a4_not_b
  PIN a5_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 132.175 238.255 147.910 238.665 ;
    END
  END a5_b
  PIN a5_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 132.770 237.475 147.900 237.930 ;
    END
  END a5_not_b
  PIN a6_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 132.175 218.285 147.910 218.695 ;
    END
  END a6_b
  PIN a6_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 132.770 217.505 147.900 217.960 ;
    END
  END a6_not_b
  PIN a7_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 132.175 198.620 147.910 199.030 ;
    END
  END a7_b
  PIN a7_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 132.770 197.840 147.900 198.295 ;
    END
  END a7_not_b
  PIN a8_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 132.215 178.780 147.950 179.190 ;
    END
  END a8_b
  PIN a8_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 132.810 178.000 147.940 178.455 ;
    END
  END a8_not_b
  PIN c0_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal3 ;
        RECT 150.720 331.265 152.465 331.575 ;
    END
  END c0_not_b
  PIN s0
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal3 ;
        RECT 148.905 328.205 150.650 328.515 ;
    END
  END s0
  PIN s0_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal3 ;
        RECT 148.935 330.250 150.680 330.560 ;
    END
  END s0_not
  PIN s1
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal3 ;
        RECT 148.775 308.475 150.520 308.785 ;
    END
  END s1
  PIN s1_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal3 ;
        RECT 148.805 310.520 150.550 310.830 ;
    END
  END s1_not
  PIN s2
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal3 ;
        RECT 148.890 288.835 150.635 289.145 ;
    END
  END s2
  PIN s2_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal3 ;
        RECT 148.920 290.880 150.665 291.190 ;
    END
  END s2_not
  PIN s3
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal3 ;
        RECT 148.890 269.035 150.635 269.345 ;
    END
  END s3
  PIN s3_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal3 ;
        RECT 148.920 271.080 150.665 271.390 ;
    END
  END s3_not
  PIN s4
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal3 ;
        RECT 148.850 249.280 150.595 249.590 ;
    END
  END s4
  PIN s4_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal3 ;
        RECT 148.880 251.325 150.625 251.635 ;
    END
  END s4_not
  PIN s5
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal3 ;
        RECT 148.890 229.565 150.635 229.875 ;
    END
  END s5
  PIN s5_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal3 ;
        RECT 148.920 231.610 150.665 231.920 ;
    END
  END s5_not
  PIN s6_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal3 ;
        RECT 148.915 211.640 150.660 211.950 ;
    END
  END s6_not
  PIN s7
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal3 ;
        RECT 148.905 189.935 150.650 190.245 ;
    END
  END s7
  PIN s7_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal3 ;
        RECT 148.935 191.980 150.680 192.290 ;
    END
  END s7_not
  PIN s6
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal3 ;
        RECT 148.885 209.595 150.630 209.905 ;
    END
  END s6
  PIN a3_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 18.135 272.830 20.595 273.135 ;
    END
  END a3_f
  PIN a3_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 18.095 272.095 20.600 272.390 ;
    END
  END a3_not_f
  PIN b3
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 18.100 271.380 20.615 271.675 ;
    END
  END b3
  PIN b3_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 18.135 270.750 20.600 271.045 ;
    END
  END b3_not
  PIN a4_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 18.005 253.120 20.465 253.425 ;
    END
  END a4_f
  PIN a4_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 17.965 252.385 20.470 252.680 ;
    END
  END a4_not_f
  PIN b4
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 17.970 251.670 20.485 251.965 ;
    END
  END b4
  PIN b4_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 18.005 251.040 20.470 251.335 ;
    END
  END b4_not
  PIN a5_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 18.135 233.360 20.595 233.665 ;
    END
  END a5_f
  PIN a5_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 18.095 232.625 20.600 232.920 ;
    END
  END a5_not_f
  PIN b5
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 18.100 231.910 20.615 232.205 ;
    END
  END b5
  PIN b5_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 18.135 231.280 20.600 231.575 ;
    END
  END b5_not
  PIN a6_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 18.085 213.550 20.545 213.855 ;
    END
  END a6_f
  PIN a6_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 18.045 212.815 20.550 213.110 ;
    END
  END a6_not_f
  PIN b6
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 18.050 212.100 20.565 212.395 ;
    END
  END b6
  PIN b6_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 18.085 211.470 20.550 211.765 ;
    END
  END b6_not
  PIN a7_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 18.055 193.755 20.515 194.060 ;
    END
  END a7_f
  PIN a7_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 18.015 193.020 20.520 193.315 ;
    END
  END a7_not_f
  PIN b7
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 18.020 192.305 20.535 192.600 ;
    END
  END b7
  PIN b7_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 18.055 191.675 20.520 191.970 ;
    END
  END b7_not
  PIN a8_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 18.205 173.960 20.665 174.265 ;
    END
  END a8_f
  PIN a8_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 18.165 173.225 20.670 173.520 ;
    END
  END a8_not_f
  PIN b8
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 18.170 172.510 20.685 172.805 ;
    END
  END b8
  PIN c0_f_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 15.050 328.050 36.160 328.345 ;
    END
  END c0_f_not
  PIN c0_f
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 15.230 328.915 35.575 329.210 ;
    END
  END c0_f
  PIN a0_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 18.185 332.070 20.645 332.375 ;
    END
  END a0_f
  PIN a0_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 18.145 331.335 20.650 331.630 ;
    END
  END a0_not_f
  PIN b0
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 18.150 330.620 20.665 330.915 ;
    END
  END b0
  PIN b0_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 18.185 329.990 20.650 330.285 ;
    END
  END b0_not
  PIN a1_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 18.140 312.380 20.600 312.685 ;
    END
  END a1_f
  PIN a1_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 18.100 311.645 20.605 311.940 ;
    END
  END a1_not_f
  PIN b1
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 18.105 310.930 20.620 311.225 ;
    END
  END b1
  PIN b1_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 18.140 310.300 20.605 310.595 ;
    END
  END b1_not
  PIN a2_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 18.330 292.670 20.790 292.975 ;
    END
  END a2_f
  PIN a2_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 18.290 291.935 20.795 292.230 ;
    END
  END a2_not_f
  PIN b2
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 18.295 291.220 20.810 291.515 ;
    END
  END b2
  PIN b2_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 18.330 290.590 20.795 290.885 ;
    END
  END b2_not
  PIN a13_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 18.115 74.515 20.620 74.810 ;
    END
  END a13_not_f
  PIN b13
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 18.120 73.800 20.635 74.095 ;
    END
  END b13
  PIN b13_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 18.155 73.170 20.620 73.465 ;
    END
  END b13_not
  PIN a14_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 18.105 55.440 20.565 55.745 ;
    END
  END a14_f
  PIN a14_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 18.065 54.705 20.570 55.000 ;
    END
  END a14_not_f
  PIN b14
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 18.070 53.990 20.585 54.285 ;
    END
  END b14
  PIN b14_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 18.105 53.360 20.570 53.655 ;
    END
  END b14_not
  PIN a15_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 18.075 35.645 20.535 35.950 ;
    END
  END a15_f
  PIN a15_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 18.035 34.910 20.540 35.205 ;
    END
  END a15_not_f
  PIN b15
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 18.040 34.195 20.555 34.490 ;
    END
  END b15
  PIN b15_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 18.075 33.565 20.540 33.860 ;
    END
  END b15_not
  PIN b8_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 18.205 171.880 20.670 172.175 ;
    END
  END b8_not
  PIN z
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 16.315 14.445 17.565 14.745 ;
    END
  END z
  PIN z_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 14.215 13.895 15.465 14.195 ;
    END
  END z_not
  PIN a9_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 18.160 154.270 20.620 154.575 ;
    END
  END a9_f
  PIN a9_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 18.120 153.535 20.625 153.830 ;
    END
  END a9_not_f
  PIN b9
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 18.125 152.820 20.640 153.115 ;
    END
  END b9
  PIN b9_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 18.160 152.190 20.625 152.485 ;
    END
  END b9_not
  PIN a10_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 18.350 134.560 20.810 134.865 ;
    END
  END a10_f
  PIN a10_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 18.310 133.825 20.815 134.120 ;
    END
  END a10_not_f
  PIN b10
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 18.315 133.110 20.830 133.405 ;
    END
  END b10
  PIN b10_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 18.350 132.480 20.815 132.775 ;
    END
  END b10_not
  PIN a11_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 18.155 114.720 20.615 115.025 ;
    END
  END a11_f
  PIN a11_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 18.115 113.985 20.620 114.280 ;
    END
  END a11_not_f
  PIN b11
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 18.120 113.270 20.635 113.565 ;
    END
  END b11
  PIN b11_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 18.155 112.640 20.620 112.935 ;
    END
  END b11_not
  PIN a12_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 18.025 95.010 20.485 95.315 ;
    END
  END a12_f
  PIN a12_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 17.985 94.275 20.490 94.570 ;
    END
  END a12_not_f
  PIN b12
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 17.990 93.560 20.505 93.855 ;
    END
  END b12
  PIN b12_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 18.025 92.930 20.490 93.225 ;
    END
  END b12_not
  PIN a13_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 18.155 75.250 20.615 75.555 ;
    END
  END a13_f
  PIN a10_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 132.170 139.410 147.905 139.820 ;
    END
  END a10_b
  PIN a10_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 132.765 138.630 147.895 139.085 ;
    END
  END a10_not_b
  PIN a11_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 132.170 119.615 147.905 120.025 ;
    END
  END a11_b
  PIN a11_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 132.765 118.835 147.895 119.290 ;
    END
  END a11_not_b
  PIN a12_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 132.090 99.860 147.825 100.270 ;
    END
  END a12_b
  PIN a12_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 132.685 99.080 147.815 99.535 ;
    END
  END a12_not_b
  PIN a13_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 132.195 80.145 147.930 80.555 ;
    END
  END a13_b
  PIN a13_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 132.790 79.365 147.920 79.820 ;
    END
  END a13_not_b
  PIN a14_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 132.195 60.175 147.930 60.585 ;
    END
  END a14_b
  PIN a14_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 132.790 59.395 147.920 59.850 ;
    END
  END a14_not_b
  PIN a15_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 132.195 40.510 147.930 40.920 ;
    END
  END a15_b
  PIN a15_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 132.790 39.730 147.920 40.185 ;
    END
  END a15_not_b
  PIN c15
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal3 ;
        RECT 103.605 11.000 111.150 11.320 ;
    END
  END c15
  PIN c15_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal3 ;
        RECT 103.620 13.430 111.140 13.750 ;
    END
  END c15_not
  PIN a9_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 132.015 159.055 147.750 159.465 ;
    END
  END a9_b
  PIN s8
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal3 ;
        RECT 148.905 170.090 150.650 170.400 ;
    END
  END s8
  PIN s8_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal3 ;
        RECT 148.935 172.135 150.680 172.445 ;
    END
  END s8_not
  PIN s9
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal3 ;
        RECT 148.805 150.365 150.550 150.675 ;
    END
  END s9
  PIN s9_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal3 ;
        RECT 148.835 152.410 150.580 152.720 ;
    END
  END s9_not
  PIN s10
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal3 ;
        RECT 148.865 130.720 150.610 131.030 ;
    END
  END s10
  PIN s10_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal3 ;
        RECT 148.895 132.765 150.640 133.075 ;
    END
  END s10_not
  PIN s11
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal3 ;
        RECT 148.865 110.930 150.610 111.240 ;
    END
  END s11
  PIN s11_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal3 ;
        RECT 148.895 112.975 150.640 113.285 ;
    END
  END s11_not
  PIN s12
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal3 ;
        RECT 148.865 91.170 150.610 91.480 ;
    END
  END s12
  PIN s12_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal3 ;
        RECT 148.895 93.215 150.640 93.525 ;
    END
  END s12_not
  PIN s13
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal3 ;
        RECT 148.890 71.460 150.635 71.770 ;
    END
  END s13
  PIN s13_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal3 ;
        RECT 148.920 73.505 150.665 73.815 ;
    END
  END s13_not
  PIN s14
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal3 ;
        RECT 148.875 51.490 150.620 51.800 ;
    END
  END s14
  PIN s14_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal3 ;
        RECT 148.905 53.535 150.650 53.845 ;
    END
  END s14_not
  PIN s15
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal3 ;
        RECT 148.900 31.825 150.645 32.135 ;
    END
  END s15
  PIN s15_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal3 ;
        RECT 148.930 33.870 150.675 34.180 ;
    END
  END s15_not
  PIN a9_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 132.610 158.275 147.740 158.730 ;
    END
  END a9_not_b
  OBS
      LAYER Nwell ;
        RECT 18.465 6.520 147.730 338.615 ;
      LAYER Metal1 ;
        RECT 9.415 6.520 156.165 338.615 ;
      LAYER Metal2 ;
        RECT 9.635 6.520 156.145 338.620 ;
      LAYER Metal3 ;
        RECT 12.115 337.600 155.440 338.570 ;
        RECT 12.115 337.370 131.895 337.600 ;
        RECT 9.560 336.590 131.895 337.370 ;
        RECT 148.230 337.370 155.440 337.600 ;
        RECT 148.230 336.590 155.770 337.370 ;
        RECT 9.560 335.810 132.490 336.590 ;
        RECT 148.220 335.810 155.770 336.590 ;
        RECT 9.560 333.285 155.770 335.810 ;
        RECT 9.560 332.675 148.980 333.285 ;
        RECT 9.560 331.930 17.885 332.675 ;
        RECT 20.945 332.375 148.980 332.675 ;
        RECT 151.515 332.375 155.770 333.285 ;
        RECT 20.945 331.930 155.770 332.375 ;
        RECT 9.560 331.035 17.845 331.930 ;
        RECT 20.950 331.875 155.770 331.930 ;
        RECT 20.950 331.215 150.420 331.875 ;
        RECT 9.560 330.320 17.850 331.035 ;
        RECT 20.965 330.965 150.420 331.215 ;
        RECT 152.765 330.965 155.770 331.875 ;
        RECT 20.965 330.860 155.770 330.965 ;
        RECT 20.965 330.320 148.635 330.860 ;
        RECT 9.560 329.690 17.885 330.320 ;
        RECT 20.950 329.950 148.635 330.320 ;
        RECT 150.980 329.950 155.770 330.860 ;
        RECT 20.950 329.690 155.770 329.950 ;
        RECT 9.560 329.510 155.770 329.690 ;
        RECT 9.560 328.645 14.930 329.510 ;
        RECT 35.875 328.815 155.770 329.510 ;
        RECT 35.875 328.645 148.605 328.815 ;
        RECT 9.560 327.750 14.750 328.645 ;
        RECT 36.460 327.905 148.605 328.645 ;
        RECT 150.950 327.905 155.770 328.815 ;
        RECT 36.460 327.750 155.770 327.905 ;
        RECT 9.560 323.895 155.770 327.750 ;
        RECT 9.560 322.395 9.975 323.895 ;
        RECT 81.545 322.395 153.695 323.895 ;
        RECT 9.560 319.125 155.770 322.395 ;
        RECT 12.120 317.875 155.445 319.125 ;
        RECT 12.120 317.625 131.695 317.875 ;
        RECT 9.560 316.865 131.695 317.625 ;
        RECT 148.030 317.625 155.445 317.875 ;
        RECT 148.030 316.865 155.770 317.625 ;
        RECT 9.560 316.085 132.290 316.865 ;
        RECT 148.020 316.085 155.770 316.865 ;
        RECT 9.560 312.985 155.770 316.085 ;
        RECT 9.560 312.240 17.840 312.985 ;
        RECT 20.900 312.240 155.770 312.985 ;
        RECT 9.560 311.345 17.800 312.240 ;
        RECT 20.905 311.525 155.770 312.240 ;
        RECT 9.560 310.630 17.805 311.345 ;
        RECT 20.920 311.130 155.770 311.525 ;
        RECT 20.920 310.630 148.505 311.130 ;
        RECT 9.560 310.000 17.840 310.630 ;
        RECT 20.905 310.220 148.505 310.630 ;
        RECT 150.850 310.220 155.770 311.130 ;
        RECT 20.905 310.000 155.770 310.220 ;
        RECT 9.560 309.085 155.770 310.000 ;
        RECT 9.560 308.175 148.475 309.085 ;
        RECT 150.820 308.175 155.770 309.085 ;
        RECT 9.560 304.125 155.770 308.175 ;
        RECT 9.560 302.625 9.975 304.125 ;
        RECT 81.545 302.625 153.695 304.125 ;
        RECT 9.560 299.485 155.770 302.625 ;
        RECT 12.110 298.230 155.435 299.485 ;
        RECT 12.110 297.985 131.850 298.230 ;
        RECT 9.560 297.220 131.850 297.985 ;
        RECT 148.185 297.985 155.435 298.230 ;
        RECT 148.185 297.220 155.770 297.985 ;
        RECT 9.560 296.440 132.445 297.220 ;
        RECT 148.175 296.440 155.770 297.220 ;
        RECT 9.560 293.275 155.770 296.440 ;
        RECT 9.560 292.530 18.030 293.275 ;
        RECT 21.090 292.530 155.770 293.275 ;
        RECT 9.560 291.635 17.990 292.530 ;
        RECT 21.095 291.815 155.770 292.530 ;
        RECT 9.560 290.920 17.995 291.635 ;
        RECT 21.110 291.490 155.770 291.815 ;
        RECT 21.110 290.920 148.620 291.490 ;
        RECT 9.560 290.290 18.030 290.920 ;
        RECT 21.095 290.580 148.620 290.920 ;
        RECT 150.965 290.580 155.770 291.490 ;
        RECT 21.095 290.290 155.770 290.580 ;
        RECT 9.560 289.445 155.770 290.290 ;
        RECT 9.560 288.535 148.590 289.445 ;
        RECT 150.935 288.535 155.770 289.445 ;
        RECT 9.560 284.430 155.770 288.535 ;
        RECT 9.560 282.930 9.975 284.430 ;
        RECT 81.545 282.930 153.695 284.430 ;
        RECT 9.560 279.690 155.770 282.930 ;
        RECT 12.120 278.435 155.445 279.690 ;
        RECT 12.120 278.190 131.850 278.435 ;
        RECT 9.560 277.425 131.850 278.190 ;
        RECT 148.185 278.190 155.445 278.435 ;
        RECT 148.185 277.425 155.770 278.190 ;
        RECT 9.560 276.645 132.445 277.425 ;
        RECT 148.175 276.645 155.770 277.425 ;
        RECT 9.560 273.435 155.770 276.645 ;
        RECT 9.560 272.690 17.835 273.435 ;
        RECT 20.895 272.690 155.770 273.435 ;
        RECT 9.560 271.795 17.795 272.690 ;
        RECT 20.900 271.975 155.770 272.690 ;
        RECT 9.560 271.080 17.800 271.795 ;
        RECT 20.915 271.690 155.770 271.975 ;
        RECT 20.915 271.080 148.620 271.690 ;
        RECT 9.560 270.450 17.835 271.080 ;
        RECT 20.900 270.780 148.620 271.080 ;
        RECT 150.965 270.780 155.770 271.690 ;
        RECT 20.900 270.450 155.770 270.780 ;
        RECT 9.560 269.645 155.770 270.450 ;
        RECT 9.560 268.735 148.590 269.645 ;
        RECT 150.935 268.735 155.770 269.645 ;
        RECT 9.560 264.695 155.770 268.735 ;
        RECT 9.560 263.195 9.975 264.695 ;
        RECT 81.545 263.195 153.695 264.695 ;
        RECT 9.560 259.940 155.770 263.195 ;
        RECT 12.130 258.680 155.455 259.940 ;
        RECT 12.130 258.440 131.770 258.680 ;
        RECT 9.560 257.670 131.770 258.440 ;
        RECT 148.105 258.440 155.455 258.680 ;
        RECT 148.105 257.670 155.770 258.440 ;
        RECT 9.560 256.890 132.365 257.670 ;
        RECT 148.095 256.890 155.770 257.670 ;
        RECT 9.560 253.725 155.770 256.890 ;
        RECT 9.560 252.980 17.705 253.725 ;
        RECT 20.765 252.980 155.770 253.725 ;
        RECT 9.560 252.085 17.665 252.980 ;
        RECT 20.770 252.265 155.770 252.980 ;
        RECT 9.560 251.370 17.670 252.085 ;
        RECT 20.785 251.935 155.770 252.265 ;
        RECT 20.785 251.370 148.580 251.935 ;
        RECT 9.560 250.740 17.705 251.370 ;
        RECT 20.770 251.025 148.580 251.370 ;
        RECT 150.925 251.025 155.770 251.935 ;
        RECT 20.770 250.740 155.770 251.025 ;
        RECT 9.560 249.890 155.770 250.740 ;
        RECT 9.560 248.980 148.550 249.890 ;
        RECT 150.895 248.980 155.770 249.890 ;
        RECT 9.560 244.940 155.770 248.980 ;
        RECT 9.560 243.440 9.975 244.940 ;
        RECT 81.545 243.440 153.695 244.940 ;
        RECT 9.560 240.230 155.770 243.440 ;
        RECT 12.095 238.965 155.420 240.230 ;
        RECT 12.095 238.730 131.875 238.965 ;
        RECT 9.560 237.955 131.875 238.730 ;
        RECT 148.210 238.730 155.420 238.965 ;
        RECT 148.210 237.955 155.770 238.730 ;
        RECT 9.560 237.175 132.470 237.955 ;
        RECT 148.200 237.175 155.770 237.955 ;
        RECT 9.560 233.965 155.770 237.175 ;
        RECT 9.560 233.220 17.835 233.965 ;
        RECT 20.895 233.220 155.770 233.965 ;
        RECT 9.560 232.325 17.795 233.220 ;
        RECT 20.900 232.505 155.770 233.220 ;
        RECT 9.560 231.610 17.800 232.325 ;
        RECT 20.915 232.220 155.770 232.505 ;
        RECT 20.915 231.610 148.620 232.220 ;
        RECT 9.560 230.980 17.835 231.610 ;
        RECT 20.900 231.310 148.620 231.610 ;
        RECT 150.965 231.310 155.770 232.220 ;
        RECT 20.900 230.980 155.770 231.310 ;
        RECT 9.560 230.175 155.770 230.980 ;
        RECT 9.560 229.265 148.590 230.175 ;
        RECT 150.935 229.265 155.770 230.175 ;
        RECT 9.560 225.190 155.770 229.265 ;
        RECT 9.560 223.690 9.995 225.190 ;
        RECT 81.565 223.690 153.715 225.190 ;
        RECT 9.560 220.265 155.770 223.690 ;
        RECT 12.130 218.995 155.455 220.265 ;
        RECT 12.130 218.765 131.875 218.995 ;
        RECT 9.560 217.985 131.875 218.765 ;
        RECT 148.210 218.765 155.455 218.995 ;
        RECT 148.210 217.985 155.770 218.765 ;
        RECT 9.560 217.205 132.470 217.985 ;
        RECT 148.200 217.205 155.770 217.985 ;
        RECT 9.560 214.155 155.770 217.205 ;
        RECT 9.560 213.410 17.785 214.155 ;
        RECT 20.845 213.410 155.770 214.155 ;
        RECT 9.560 212.515 17.745 213.410 ;
        RECT 20.850 212.695 155.770 213.410 ;
        RECT 9.560 211.800 17.750 212.515 ;
        RECT 20.865 212.250 155.770 212.695 ;
        RECT 20.865 211.800 148.615 212.250 ;
        RECT 9.560 211.170 17.785 211.800 ;
        RECT 20.850 211.340 148.615 211.800 ;
        RECT 150.960 211.340 155.770 212.250 ;
        RECT 20.850 211.170 155.770 211.340 ;
        RECT 9.560 210.205 155.770 211.170 ;
        RECT 9.560 209.295 148.585 210.205 ;
        RECT 150.930 209.295 155.770 210.205 ;
        RECT 9.560 205.245 155.770 209.295 ;
        RECT 9.560 203.745 9.995 205.245 ;
        RECT 81.565 203.745 153.715 205.245 ;
        RECT 9.560 200.580 155.770 203.745 ;
        RECT 12.110 199.330 155.435 200.580 ;
        RECT 12.110 199.080 131.875 199.330 ;
        RECT 9.560 198.320 131.875 199.080 ;
        RECT 148.210 199.080 155.435 199.330 ;
        RECT 148.210 198.320 155.770 199.080 ;
        RECT 9.560 197.540 132.470 198.320 ;
        RECT 148.200 197.540 155.770 198.320 ;
        RECT 9.560 194.360 155.770 197.540 ;
        RECT 9.560 193.615 17.755 194.360 ;
        RECT 20.815 193.615 155.770 194.360 ;
        RECT 9.560 192.720 17.715 193.615 ;
        RECT 20.820 192.900 155.770 193.615 ;
        RECT 9.560 192.005 17.720 192.720 ;
        RECT 20.835 192.590 155.770 192.900 ;
        RECT 20.835 192.005 148.635 192.590 ;
        RECT 9.560 191.375 17.755 192.005 ;
        RECT 20.820 191.680 148.635 192.005 ;
        RECT 150.980 191.680 155.770 192.590 ;
        RECT 20.820 191.375 155.770 191.680 ;
        RECT 9.560 190.545 155.770 191.375 ;
        RECT 9.560 189.635 148.605 190.545 ;
        RECT 150.950 189.635 155.770 190.545 ;
        RECT 9.560 185.550 155.770 189.635 ;
        RECT 9.560 184.050 9.975 185.550 ;
        RECT 81.545 184.050 153.695 185.550 ;
        RECT 9.560 180.740 155.770 184.050 ;
        RECT 12.110 179.490 155.435 180.740 ;
        RECT 12.110 179.240 131.915 179.490 ;
        RECT 9.560 178.480 131.915 179.240 ;
        RECT 148.250 179.240 155.435 179.490 ;
        RECT 148.250 178.480 155.770 179.240 ;
        RECT 9.560 177.700 132.510 178.480 ;
        RECT 148.240 177.700 155.770 178.480 ;
        RECT 9.560 174.565 155.770 177.700 ;
        RECT 9.560 173.820 17.905 174.565 ;
        RECT 20.965 173.820 155.770 174.565 ;
        RECT 9.560 172.925 17.865 173.820 ;
        RECT 20.970 173.105 155.770 173.820 ;
        RECT 9.560 172.210 17.870 172.925 ;
        RECT 20.985 172.745 155.770 173.105 ;
        RECT 20.985 172.210 148.635 172.745 ;
        RECT 9.560 171.580 17.905 172.210 ;
        RECT 20.970 171.835 148.635 172.210 ;
        RECT 150.980 171.835 155.770 172.745 ;
        RECT 20.970 171.580 155.770 171.835 ;
        RECT 9.560 170.700 155.770 171.580 ;
        RECT 9.560 169.790 148.605 170.700 ;
        RECT 150.950 169.790 155.770 170.700 ;
        RECT 9.560 165.780 155.770 169.790 ;
        RECT 9.560 164.280 10.030 165.780 ;
        RECT 81.600 164.280 153.750 165.780 ;
        RECT 9.560 161.045 155.770 164.280 ;
        RECT 12.120 159.765 155.445 161.045 ;
        RECT 12.120 159.545 131.715 159.765 ;
        RECT 9.560 158.755 131.715 159.545 ;
        RECT 148.050 159.545 155.445 159.765 ;
        RECT 148.050 158.755 155.770 159.545 ;
        RECT 9.560 157.975 132.310 158.755 ;
        RECT 148.040 157.975 155.770 158.755 ;
        RECT 9.560 154.875 155.770 157.975 ;
        RECT 9.560 154.130 17.860 154.875 ;
        RECT 20.920 154.130 155.770 154.875 ;
        RECT 9.560 153.235 17.820 154.130 ;
        RECT 20.925 153.415 155.770 154.130 ;
        RECT 9.560 152.520 17.825 153.235 ;
        RECT 20.940 153.020 155.770 153.415 ;
        RECT 20.940 152.520 148.535 153.020 ;
        RECT 9.560 151.890 17.860 152.520 ;
        RECT 20.925 152.110 148.535 152.520 ;
        RECT 150.880 152.110 155.770 153.020 ;
        RECT 20.925 151.890 155.770 152.110 ;
        RECT 9.560 150.975 155.770 151.890 ;
        RECT 9.560 150.065 148.505 150.975 ;
        RECT 150.850 150.065 155.770 150.975 ;
        RECT 9.560 146.045 155.770 150.065 ;
        RECT 9.560 144.545 9.975 146.045 ;
        RECT 81.545 144.545 153.695 146.045 ;
        RECT 9.560 141.380 155.770 144.545 ;
        RECT 12.120 140.120 155.445 141.380 ;
        RECT 12.120 139.880 131.870 140.120 ;
        RECT 9.560 139.110 131.870 139.880 ;
        RECT 148.205 139.880 155.445 140.120 ;
        RECT 148.205 139.110 155.770 139.880 ;
        RECT 9.560 138.330 132.465 139.110 ;
        RECT 148.195 138.330 155.770 139.110 ;
        RECT 9.560 135.165 155.770 138.330 ;
        RECT 9.560 134.420 18.050 135.165 ;
        RECT 21.110 134.420 155.770 135.165 ;
        RECT 9.560 133.525 18.010 134.420 ;
        RECT 21.115 133.705 155.770 134.420 ;
        RECT 9.560 132.810 18.015 133.525 ;
        RECT 21.130 133.375 155.770 133.705 ;
        RECT 21.130 132.810 148.595 133.375 ;
        RECT 9.560 132.180 18.050 132.810 ;
        RECT 21.115 132.465 148.595 132.810 ;
        RECT 150.940 132.465 155.770 133.375 ;
        RECT 21.115 132.180 155.770 132.465 ;
        RECT 9.560 131.330 155.770 132.180 ;
        RECT 9.560 130.420 148.565 131.330 ;
        RECT 150.910 130.420 155.770 131.330 ;
        RECT 9.560 126.365 155.770 130.420 ;
        RECT 9.560 124.865 9.975 126.365 ;
        RECT 81.545 124.865 153.695 126.365 ;
        RECT 9.560 121.540 155.770 124.865 ;
        RECT 12.110 120.325 155.435 121.540 ;
        RECT 12.110 120.040 131.870 120.325 ;
        RECT 9.560 119.315 131.870 120.040 ;
        RECT 148.205 120.040 155.435 120.325 ;
        RECT 148.205 119.315 155.770 120.040 ;
        RECT 9.560 118.535 132.465 119.315 ;
        RECT 148.195 118.535 155.770 119.315 ;
        RECT 9.560 115.325 155.770 118.535 ;
        RECT 9.560 114.580 17.855 115.325 ;
        RECT 20.915 114.580 155.770 115.325 ;
        RECT 9.560 113.685 17.815 114.580 ;
        RECT 20.920 113.865 155.770 114.580 ;
        RECT 9.560 112.970 17.820 113.685 ;
        RECT 20.935 113.585 155.770 113.865 ;
        RECT 20.935 112.970 148.595 113.585 ;
        RECT 9.560 112.340 17.855 112.970 ;
        RECT 20.920 112.675 148.595 112.970 ;
        RECT 150.940 112.675 155.770 113.585 ;
        RECT 20.920 112.340 155.770 112.675 ;
        RECT 9.560 111.540 155.770 112.340 ;
        RECT 9.560 110.630 148.565 111.540 ;
        RECT 150.910 110.630 155.770 111.540 ;
        RECT 9.560 106.575 155.770 110.630 ;
        RECT 9.560 105.075 9.995 106.575 ;
        RECT 81.565 105.075 153.715 106.575 ;
        RECT 9.560 101.850 155.770 105.075 ;
        RECT 12.110 100.570 155.435 101.850 ;
        RECT 12.110 100.350 131.790 100.570 ;
        RECT 9.560 99.560 131.790 100.350 ;
        RECT 148.125 100.350 155.435 100.570 ;
        RECT 148.125 99.560 155.770 100.350 ;
        RECT 9.560 98.780 132.385 99.560 ;
        RECT 148.115 98.780 155.770 99.560 ;
        RECT 9.560 95.615 155.770 98.780 ;
        RECT 9.560 94.870 17.725 95.615 ;
        RECT 20.785 94.870 155.770 95.615 ;
        RECT 9.560 93.975 17.685 94.870 ;
        RECT 20.790 94.155 155.770 94.870 ;
        RECT 9.560 93.260 17.690 93.975 ;
        RECT 20.805 93.825 155.770 94.155 ;
        RECT 20.805 93.260 148.595 93.825 ;
        RECT 9.560 92.630 17.725 93.260 ;
        RECT 20.790 92.915 148.595 93.260 ;
        RECT 150.940 92.915 155.770 93.825 ;
        RECT 20.790 92.630 155.770 92.915 ;
        RECT 9.560 91.780 155.770 92.630 ;
        RECT 9.560 90.870 148.565 91.780 ;
        RECT 150.910 90.870 155.770 91.780 ;
        RECT 9.560 86.795 155.770 90.870 ;
        RECT 9.560 85.295 10.010 86.795 ;
        RECT 81.580 85.295 153.730 86.795 ;
        RECT 9.560 82.110 155.770 85.295 ;
        RECT 12.110 80.855 155.435 82.110 ;
        RECT 12.110 80.610 131.895 80.855 ;
        RECT 9.560 79.845 131.895 80.610 ;
        RECT 148.230 80.610 155.435 80.855 ;
        RECT 148.230 79.845 155.770 80.610 ;
        RECT 9.560 79.065 132.490 79.845 ;
        RECT 148.220 79.065 155.770 79.845 ;
        RECT 9.560 75.855 155.770 79.065 ;
        RECT 9.560 75.110 17.855 75.855 ;
        RECT 20.915 75.110 155.770 75.855 ;
        RECT 9.560 74.215 17.815 75.110 ;
        RECT 20.920 74.395 155.770 75.110 ;
        RECT 9.560 73.500 17.820 74.215 ;
        RECT 20.935 74.115 155.770 74.395 ;
        RECT 20.935 73.500 148.620 74.115 ;
        RECT 9.560 72.870 17.855 73.500 ;
        RECT 20.920 73.205 148.620 73.500 ;
        RECT 150.965 73.205 155.770 74.115 ;
        RECT 20.920 72.870 155.770 73.205 ;
        RECT 9.560 72.070 155.770 72.870 ;
        RECT 9.560 71.160 148.590 72.070 ;
        RECT 150.935 71.160 155.770 72.070 ;
        RECT 9.560 67.065 155.770 71.160 ;
        RECT 9.560 65.565 9.915 67.065 ;
        RECT 81.485 65.565 153.635 67.065 ;
        RECT 9.560 62.180 155.770 65.565 ;
        RECT 12.145 60.885 155.470 62.180 ;
        RECT 12.145 60.680 131.895 60.885 ;
        RECT 9.560 59.875 131.895 60.680 ;
        RECT 148.230 60.680 155.470 60.885 ;
        RECT 148.230 59.875 155.770 60.680 ;
        RECT 9.560 59.095 132.490 59.875 ;
        RECT 148.220 59.095 155.770 59.875 ;
        RECT 9.560 56.045 155.770 59.095 ;
        RECT 9.560 55.300 17.805 56.045 ;
        RECT 20.865 55.300 155.770 56.045 ;
        RECT 9.560 54.405 17.765 55.300 ;
        RECT 20.870 54.585 155.770 55.300 ;
        RECT 9.560 53.690 17.770 54.405 ;
        RECT 20.885 54.145 155.770 54.585 ;
        RECT 20.885 53.690 148.605 54.145 ;
        RECT 9.560 53.060 17.805 53.690 ;
        RECT 20.870 53.235 148.605 53.690 ;
        RECT 150.950 53.235 155.770 54.145 ;
        RECT 20.870 53.060 155.770 53.235 ;
        RECT 9.560 52.100 155.770 53.060 ;
        RECT 9.560 51.190 148.575 52.100 ;
        RECT 150.920 51.190 155.770 52.100 ;
        RECT 9.560 47.110 155.770 51.190 ;
        RECT 9.560 45.610 10.010 47.110 ;
        RECT 81.580 45.610 153.730 47.110 ;
        RECT 9.560 42.540 155.770 45.610 ;
        RECT 12.125 41.220 155.450 42.540 ;
        RECT 12.125 41.040 131.895 41.220 ;
        RECT 9.560 40.210 131.895 41.040 ;
        RECT 148.230 41.040 155.450 41.220 ;
        RECT 148.230 40.210 155.770 41.040 ;
        RECT 9.560 39.430 132.490 40.210 ;
        RECT 148.220 39.430 155.770 40.210 ;
        RECT 9.560 36.250 155.770 39.430 ;
        RECT 9.560 35.505 17.775 36.250 ;
        RECT 20.835 35.505 155.770 36.250 ;
        RECT 9.560 34.610 17.735 35.505 ;
        RECT 20.840 34.790 155.770 35.505 ;
        RECT 9.560 33.895 17.740 34.610 ;
        RECT 20.855 34.480 155.770 34.790 ;
        RECT 20.855 33.895 148.630 34.480 ;
        RECT 9.560 33.265 17.775 33.895 ;
        RECT 20.840 33.570 148.630 33.895 ;
        RECT 150.975 33.570 155.770 34.480 ;
        RECT 20.840 33.265 155.770 33.570 ;
        RECT 9.560 32.435 155.770 33.265 ;
        RECT 9.560 31.525 148.600 32.435 ;
        RECT 150.945 31.525 155.770 32.435 ;
        RECT 9.560 27.485 155.770 31.525 ;
        RECT 9.560 25.985 10.025 27.485 ;
        RECT 81.595 25.985 153.745 27.485 ;
        RECT 9.560 22.760 155.770 25.985 ;
        RECT 12.110 21.260 155.435 22.760 ;
        RECT 9.560 15.045 155.770 21.260 ;
        RECT 9.560 14.495 16.015 15.045 ;
        RECT 9.560 13.595 13.915 14.495 ;
        RECT 15.765 14.145 16.015 14.495 ;
        RECT 17.865 14.145 155.770 15.045 ;
        RECT 15.765 14.050 155.770 14.145 ;
        RECT 15.765 13.595 103.320 14.050 ;
        RECT 9.560 13.130 103.320 13.595 ;
        RECT 111.440 13.130 155.770 14.050 ;
        RECT 9.560 11.620 155.770 13.130 ;
        RECT 9.560 10.700 103.305 11.620 ;
        RECT 111.450 10.700 155.770 11.620 ;
        RECT 9.560 7.710 155.770 10.700 ;
        RECT 9.560 6.510 9.990 7.710 ;
        RECT 81.560 6.510 153.710 7.710 ;
  END
END 16b_FA
END LIBRARY

