`default_nettype none

(* blackbox *)
module CCNOT (
    inout wire VDD,
    inout wire VSS,
    inout wire a,
    inout wire a_not,
    inout wire b,
    inout wire b_not,
    inout wire c,
    inout wire c_not,
    inout wire r_not,
    inout wire r,
    inout wire p,
    inout wire p_not,
    inout wire q,
    inout wire q_not,
);

endmodule

