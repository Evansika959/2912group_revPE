* Extracted by KLayout with GF180MCU LVS runset on : 03/12/2025 14:02

.SUBCKT 8b_mult b6_c5 vss x0_b0_f x1_b0_f x2_b0_f x3_b0_f x4_b0_f x5_b0_f
+ x6_b0_f p15_not x0_b0_f_not x1_b0_f_not x2_b0_f_not x3_b0_f_not x4_b0_f_not
+ x5_b0_f_not x6_b0_f_not p15 vdd
+ a7_not|b0_p7_not|b1_p7_not|b2_p7_not|b4_p7_not|b5_p7_not|b6_p7_not|b7_p7_not
+ a7|b0_p7|b1_p7|b2_p7|b3_p7|b4_p7|b5_p7|b6_p7|b7_p7 b2_p7_not|b3_p7_not
+ b1_c7_not x0_a7_b_not x0_a7_b b2_c7_not b2_r7_b_not b2_r7_b b3_c7_not
+ b3_r7_b_not b3_r7_b b4_c7_not b4_r7_b_not b4_r7_b b5_c7_not b5_r7_b_not
+ b5_r7_b b6_c7_not b6_r7_b_not b6_r7_b p14 p14_not
+ b1_not|b1_q0_not|b1_q1_not|b1_q2_not|b1_q3_not|b1_q4_not|b1_q5_not|b1_q6_not|b1_q7_not
+ b2_not|b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not
+ b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b3_not|b3_q0_not|b3_q1_not|b3_q2_not|b3_q3_not|b3_q4_not|b3_q5_not|b3_q6_not|b3_q7_not
+ b2_q0_not|b2_q1_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b4_not|b4_q7_not
+ b5_not|b5_q0_not|b5_q1_not|b5_q2_not|b5_q3_not|b5_q4_not|b5_q5_not|b5_q6_not|b5_q7_not
+ b6_not|b6_q0_not|b6_q1_not|b6_q2_not|b6_q3_not|b6_q4_not|b6_q5_not|b6_q6_not|b6_q7_not
+ b7_not|b7_q0_not|b7_q1_not|b7_q2_not|b7_q3_not|b7_q4_not|b7_q5_not|b7_q6_not|b7_q7_not
+ b1_c7 b1|b1_q0|b1_q1|b1_q2|b1_q3|b1_q4|b1_q5|b1_q6|b1_q7
+ b2|b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7 b2_c7
+ b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b3|b3_q0|b3_q1|b3_q2|b3_q3|b3_q4|b3_q5|b3_q6|b3_q7
+ b3_c7 b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b4|b4_q7 b4_c7
+ b5|b5_q0|b5_q1|b5_q2|b5_q3|b5_q4|b5_q5|b5_q6|b5_q7 b5_c7
+ b6|b6_q0|b6_q1|b6_q2|b6_q3|b6_q4|b6_q5|b6_q6|b6_q7 b6_c7
+ b1_q3|b7|b7_q0|b7_q1|b7_q2|b7_q4|b7_q5|b7_q6|b7_q7 x0_a7_f x0_a7_f_not
+ a6_not|b0_p6_not|b1_p6_not|b3_p6_not|b4_p6_not|b5_p6_not|b6_p6_not|b7_p6_not
+ a6|b0_p6|b1_p6|b3_p6|b4_p6|b5_p6|b6_p6|b7_p6 b1_c6_not b1_c6 b0_c7_not b0_c7
+ b0_r7_b_not b0_r7_b b2_c6_not b2_r6_b_not b2_r6_b b3_c6_not b3_r6_b_not
+ b3_r6_b b4_c6_not b4_r6_b_not b4_r6_b b5_c6_not b5_r6_b_not b5_r6_b b6_c6_not
+ b6_r6_b_not b6_r6_b p13 p13_not
+ b0_not|b0_q0_not|b0_q1_not|b0_q3_not|b0_q4_not|b0_q5_not|b0_q6_not|b0_q7_not|b1_q2_not
+ b0|b0_q0|b0_q1|b0_q2|b0_q3|b0_q4|b0_q5|b0_q6|b0_q7 b2_c6 b3_c6 b4_c6 b5_c6
+ b6_c6
+ a5_not|b0_p5_not|b1_p5_not|b2_p5_not|b3_p5_not|b5_p5_not|b6_p5_not|b7_p5_not
+ a5|b0_p5|b1_p5|b3_p5|b4_p5|b5_p5|b6_p5|b7_p5 b1_c5_not b0_c6_not b0_r6_b_not
+ b0_r6_b b2_c5_not b2_r5_b_not b2_r5_b b3_r5_b_not b3_r5_b b4_r5_b_not b4_r5_b
+ b5_r5_b_not b5_r5_b b6_c5_not b6_r5_b_not b6_r5_b p12_not b1_c5 b0_c6 p12
+ b2_c5 b3_c5 b5_c5
+ a4_not|b0_p4_not|b1_p4_not|b2_p4_not|b3_p4_not|b5_p4_not|b6_p4_not|b7_p4_not
+ a4|b0_p4|b1_p4|b2_p4|b3_p4|b4_p4|b5_p4|b6_p4|b7_p4 b1_c4_not b0_c5_not
+ b0_r5_b_not b0_r5_b b2_c4_not b2_r4_b_not b2_r4_b b3_r4_b_not b3_r4_b
+ b4_r4_b_not b4_r4_b b5_r4_b_not b5_r4_b b6_c4_not b6_r4_b_not b6_r4_b p11
+ p11_not b1_c4 b0_c5 b6_c4 b2_c4
+ a3_not|b0_p3_not|b1_p3_not|b2_p3_not|b3_p3_not|b5_p3_not|b6_p3_not|b7_p3_not
+ a3|b0_p3|b1_p3|b2_p3|b3_p3|b5_p3|b6_p3|b7_p3 b1_c3_not b0_c4_not b0_r4_b_not
+ b0_r4_b b2_c2_not b2_r3_b_not b2_r3_b b3_c2_not b3_r3_b_not b3_r3_b b4_c2_not
+ b4_r3_b_not b4_r3_b b5_c2_not b5_r3_b_not b5_r3_b b6_c2_not|b6_c3_not
+ b6_r3_b_not b6_r3_b b6_c2_not p10 p10_not b1_c3 b0_c4 b2_c2 b3_c2 b4_c2 b5_c2
+ b6_c2 b6_c2|b6_c3
+ a2_not|b0_p2_not|b1_p2_not|b2_p2_not|b3_p2_not|b5_p2_not|b6_p2_not|b7_p2_not
+ a2|b0_p2|b1_p2|b2_p2|b3_p2|b4_p2|b5_p2|b6_p2|b7_p2 b1_c2_not b0_c3_not
+ b2_r2_b_not b2_r2_b b3_r2_b_not b3_r2_b b4_r2_b_not b4_r2_b b5_r2_b_not
+ b5_r2_b b6_r2_b_not b6_r2_b p9 p9_not b1_c2 b0_c3
+ a1_not|b0_p1_not|b1_p1_not|b2_p1_not|b3_p1_not|b4_p1_not|b5_p1_not|b6_p1_not|b7_p1_not
+ b1_c1_not a1|b0_p1|b1_p1|b2_p1|b3_p1|b4_p1|b5_p1|b6_p1|b7_p1 b2_r1_b_not
+ b2_r1_b b2_c1_not b3_r1_b_not b3_r1_b b4_r1_b_not b4_r1_b b5_r1_b_not b5_r1_b
+ b6_r1_b_not b6_r1_b b0_c2_not b6_c1_not p8 p8_not b1_c1 b0_c2 b2_c1 b3_c1
+ b4_c1 b5_c1 b6_c1
+ a0_not|b0_p0_not|b1_p0_not|b2_p0_not|b3_p0_not|b5_p0_not|b6_p0_not|b7_p0_not
+ a0|b0_p0|b1_p0|b2_p0|b3_p0|b4_p0|b5_p0|b6_p0|b7_p0 b1_c0_not b0_c1_not
+ b2_c0_not b2_r0_b_not b2_r0_b b3_r0_b_not b3_r0_b b4_r0_b_not b4_r0_b
+ b5_r0_b_not b5_r0_b b6_c0_not b6_r0_b_not b6_r0_b x0_c0_b x0_c0_b_not p1
+ p1_not p2 p2_not p3 p3_not p4 p4_not p5 p5_not p6 p6_not p7 p7_not b1_c0
+ b0_c1 b2_c0 x0_c0_f x0_c0_f_not b6_c0 b0_c0_not p0_not b0_c0 p0
M$1 x2_b0_f_not \$166 \$17 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$2 \$15 \$80 x2_b0_f_not vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$3 x2_b0_f \$166 \$15 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$4 x3_b0_f_not \$173 \$19 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$5 x4_b0_f_not \$180 \$21 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$6 x5_b0_f_not \$187 \$23 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$7 x6_b0_f_not \$194 p15_not vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$8 x0_b0_f_not \$152 \$28 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$9 x1_b0_f_not \$159 \$31 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$10 \$34 \$82 x3_b0_f_not vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$11 x3_b0_f \$173 \$34 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$12 \$36 \$84 x4_b0_f_not vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$13 x4_b0_f \$180 \$36 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$14 \$38 \$86 x5_b0_f_not vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$15 x5_b0_f \$187 \$38 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$16 p15 \$88 x6_b0_f_not vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$17 x6_b0_f \$194 p15 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$18 \$27 \$76 x0_b0_f_not vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$19 x0_b0_f \$152 \$27 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$20 \$28 \$76 x0_b0_f vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P AD=0.60515P
+ PS=3.52U PD=3.45U
M$21 \$30 \$78 x1_b0_f_not vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$22 x1_b0_f \$159 \$30 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$23 \$31 \$78 x1_b0_f vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P AD=0.60515P
+ PS=3.52U PD=3.45U
M$24 \$30 \$165 \$289 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$25 \$223 \$165 \$145 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$26 \$17 \$80 x2_b0_f vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P AD=0.60515P
+ PS=3.52U PD=3.45U
M$27 \$290 b3_r7_b_not \$145 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$28 \$145 b3_r7_b \$291 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$29 \$292 \$291 \$289 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$30 \$289 \$290 \$293 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$31 \$19 \$82 x3_b0_f vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P AD=0.60515P
+ PS=3.52U PD=3.45U
M$32 \$21 \$84 x4_b0_f vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P AD=0.60515P
+ PS=3.52U PD=3.45U
M$33 \$23 \$86 x5_b0_f vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P AD=0.60515P
+ PS=3.52U PD=3.45U
M$34 p15_not \$88 x6_b0_f vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$35 \$287 \$163 \$30 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$36 \$31 \$165 \$287 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$37 \$288 \$163 \$223 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$38 \$451 \$165 \$288 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$39 \$288 b3_r7_b \$290 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$40 \$287 \$290 \$292 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$41 \$298 b4_r7_b_not \$146 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$42 \$146 b4_r7_b \$299 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$43 \$300 \$299 \$296 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$44 \$296 \$298 \$301 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$45 \$306 b5_r7_b_not \$147 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$46 \$147 b5_r7_b \$307 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$47 \$308 \$307 \$304 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$48 \$304 \$306 \$309 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$49 \$314 b6_r7_b_not \$148 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$50 \$148 b6_r7_b \$315 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$51 \$316 \$315 \$312 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$52 \$312 \$314 \$317 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$53 \$322 \$195 \$149 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$54 \$149 \$196 \$323 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$55 p14 \$323 \$320 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$56 \$320 \$322 p14_not vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$57 \$142 x0_a7_b \$275 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$58 \$272 \$274 \$277 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$59 \$143 b2_r7_b \$283 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$60 \$280 \$282 \$285 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$61 \$295 \$170 \$15 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$62 \$15 \$172 \$296 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$63 \$297 \$170 \$224 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$64 \$224 \$172 \$146 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$65 \$297 b4_r7_b \$298 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$66 \$295 \$298 \$300 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$67 \$303 \$177 \$34 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$68 \$34 \$179 \$304 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$69 \$305 \$177 \$225 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$70 \$225 \$179 \$147 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$71 \$305 b5_r7_b \$306 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$72 \$303 \$306 \$308 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$73 \$311 \$184 \$36 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$74 \$36 \$186 \$312 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$75 \$313 \$184 \$226 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$76 \$226 \$186 \$148 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$77 \$313 b6_r7_b \$314 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$78 \$311 \$314 \$316 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$79 \$319 \$191 \$38 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$80 \$38 \$193 \$320 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$81 \$321 \$191 \$227 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$82 \$227 \$193 \$149 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$83 \$321 \$196 \$322 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$84 \$319 \$322 p14 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$85 \$271 x0_a7_f_not \$220 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$86 \$151 x0_a7_f \$271 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$87 \$272 x0_a7_f_not \$151 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$88 \$220 x0_a7_f \$272 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$89 \$273 x0_a7_f_not \$221 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$90 \$608 x0_a7_f \$273 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$91 \$142 x0_a7_f_not \$608 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$92 \$221 x0_a7_f \$142 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$93 \$274 x0_a7_b_not \$142 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$94 \$273 x0_a7_b \$274 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$95 \$275 x0_a7_b_not \$273 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$96 \$276 \$275 \$272 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$97 \$271 \$274 \$276 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$98 \$277 \$275 \$271 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P AD=0.60515P
+ PS=3.52U PD=3.45U
M$99 \$279 \$156 \$27 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$100 \$28 \$158 \$279 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$101 \$280 \$156 \$28 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P AD=0.60515P
+ PS=3.52U PD=3.45U
M$102 \$27 \$158 \$280 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$103 \$281 \$156 \$222 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$104 \$613 \$158 \$281 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$105 \$143 \$156 \$613 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P AD=0.60515P
+ PS=3.52U PD=3.45U
M$106 \$222 \$158 \$143 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$107 \$282 b2_r7_b_not \$143 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$108 \$281 b2_r7_b \$282 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$109 \$283 b2_r7_b_not \$281 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$110 \$284 \$283 \$280 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$111 \$279 \$282 \$284 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$112 \$285 \$283 \$279 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P AD=0.60515P
+ PS=3.52U PD=3.45U
M$113 \$289 \$163 \$31 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P AD=0.60515P
+ PS=3.52U PD=3.45U
M$114 \$145 \$163 \$451 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P AD=0.60515P
+ PS=3.52U PD=3.45U
M$115 \$291 b3_r7_b_not \$288 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$116 \$293 \$291 \$287 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P AD=0.60515P
+ PS=3.52U PD=3.45U
M$117 \$17 \$172 \$295 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$118 \$296 \$170 \$17 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P AD=0.60515P
+ PS=3.52U PD=3.45U
M$119 \$622 \$172 \$297 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$120 \$146 \$170 \$622 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P AD=0.60515P
+ PS=3.52U PD=3.45U
M$121 \$299 b4_r7_b_not \$297 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$122 \$301 \$299 \$295 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P AD=0.60515P
+ PS=3.52U PD=3.45U
M$123 \$19 \$179 \$303 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$124 \$304 \$177 \$19 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P AD=0.60515P
+ PS=3.52U PD=3.45U
M$125 \$627 \$179 \$305 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$126 \$147 \$177 \$627 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P AD=0.60515P
+ PS=3.52U PD=3.45U
M$127 \$307 b5_r7_b_not \$305 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$128 \$309 \$307 \$303 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P AD=0.60515P
+ PS=3.52U PD=3.45U
M$129 \$21 \$186 \$311 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$130 \$312 \$184 \$21 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P AD=0.60515P
+ PS=3.52U PD=3.45U
M$131 \$632 \$186 \$313 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$132 \$148 \$184 \$632 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P AD=0.60515P
+ PS=3.52U PD=3.45U
M$133 \$315 b6_r7_b_not \$313 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$134 \$317 \$315 \$311 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P AD=0.60515P
+ PS=3.52U PD=3.45U
M$135 \$23 \$193 \$319 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$136 \$320 \$191 \$23 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P AD=0.60515P
+ PS=3.52U PD=3.45U
M$137 \$637 \$193 \$321 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$138 \$149 \$191 \$637 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P AD=0.60515P
+ PS=3.52U PD=3.45U
M$139 \$323 \$195 \$321 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P AD=0.60515P
+ PS=3.52U PD=3.45U
M$140 p14_not \$323 \$319 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$141 \$220 b1|b1_q0|b1_q1|b1_q2|b1_q3|b1_q4|b1_q5|b1_q6|b1_q7 b1_c7_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$142 \$683
+ b1_not|b1_q0_not|b1_q1_not|b1_q2_not|b1_q3_not|b1_q4_not|b1_q5_not|b1_q6_not|b1_q7_not
+ \$220 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$143 b1_c7
+ a7_not|b0_p7_not|b1_p7_not|b2_p7_not|b4_p7_not|b5_p7_not|b6_p7_not|b7_p7_not
+ \$683 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$144 \$684
+ a7_not|b0_p7_not|b1_p7_not|b2_p7_not|b4_p7_not|b5_p7_not|b6_p7_not|b7_p7_not
+ b1_c7_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$145 \$151
+ b1_not|b1_q0_not|b1_q1_not|b1_q2_not|b1_q3_not|b1_q4_not|b1_q5_not|b1_q6_not|b1_q7_not
+ \$684 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$146 b1_c7 b1|b1_q0|b1_q1|b1_q2|b1_q3|b1_q4|b1_q5|b1_q6|b1_q7 \$151 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$147 \$76 \$271 x0_a7_f_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$148 \$685 \$272 \$76 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$149 x0_a7_f \$142 \$685 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$150 \$686 \$142 x0_a7_f_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$151 \$152 \$272 \$686 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$152 x0_a7_f \$271 \$152 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$153 x0_a7_b_not \$271 \$76 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$154 \$687 \$272 x0_a7_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$155 \$152 \$142 \$687 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$156 \$688 \$142 \$76 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$157 x0_a7_b \$272 \$688 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$158 \$152 \$271 x0_a7_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$159 \$156 b2|b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7 b2_c7_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$160 \$689
+ b2_not|b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not
+ \$156 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$161 b2_c7
+ a7_not|b0_p7_not|b1_p7_not|b2_p7_not|b4_p7_not|b5_p7_not|b6_p7_not|b7_p7_not
+ \$689 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$162 \$690
+ a7_not|b0_p7_not|b1_p7_not|b2_p7_not|b4_p7_not|b5_p7_not|b6_p7_not|b7_p7_not
+ b2_c7_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$163 \$158
+ b2_not|b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not
+ \$690 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$164 b2_c7 b2|b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7 \$158 vdd pfet_03v3
+ L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$165 \$78 \$279 \$156 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$166 \$691 \$280 \$78 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$167 \$158 \$143 \$691 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$168 \$692 \$143 \$156 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$169 \$159 \$280 \$692 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$170 \$158 \$279 \$159 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$171 b2_r7_b_not \$279 \$78 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$172 \$693 \$280 b2_r7_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$173 \$159 \$143 \$693 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$174 \$694 \$143 \$78 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$175 b2_r7_b \$280 \$694 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$176 \$159 \$279 b2_r7_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$177 \$163
+ b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b3|b3_q0|b3_q1|b3_q2|b3_q3|b3_q4|b3_q5|b3_q6|b3_q7
+ b3_c7_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$178 \$695
+ b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b3_not|b3_q0_not|b3_q1_not|b3_q2_not|b3_q3_not|b3_q4_not|b3_q5_not|b3_q6_not|b3_q7_not
+ \$163 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$179 b3_c7 b2_p7_not|b3_p7_not \$695 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$180 \$696 b2_p7_not|b3_p7_not b3_c7_not vdd pfet_03v3 L=0.28U W=0.42U
+ AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$181 \$165
+ b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b3_not|b3_q0_not|b3_q1_not|b3_q2_not|b3_q3_not|b3_q4_not|b3_q5_not|b3_q6_not|b3_q7_not
+ \$696 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$182 b3_c7
+ b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b3|b3_q0|b3_q1|b3_q2|b3_q3|b3_q4|b3_q5|b3_q6|b3_q7
+ \$165 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$183 \$80 \$287 \$163 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$184 \$697 \$289 \$80 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$185 \$165 \$145 \$697 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$186 \$698 \$145 \$163 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$187 \$166 \$289 \$698 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$188 \$165 \$287 \$166 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$189 b3_r7_b_not \$287 \$80 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$190 \$699 \$289 b3_r7_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$191 \$166 \$145 \$699 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$192 \$700 \$145 \$80 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$193 b3_r7_b \$289 \$700 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$194 \$166 \$287 b3_r7_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$195 \$82 \$295 \$170 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$196 \$701 \$296 \$82 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$197 \$172 \$146 \$701 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$198 \$702 \$146 \$170 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$199 \$173 \$296 \$702 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$200 \$172 \$295 \$173 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$201 b4_r7_b_not \$295 \$82 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$202 \$703 \$296 b4_r7_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$203 \$173 \$146 \$703 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$204 \$704 \$146 \$82 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$205 b4_r7_b \$296 \$704 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$206 \$173 \$295 b4_r7_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$207 \$84 \$303 \$177 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$208 \$705 \$304 \$84 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$209 \$179 \$147 \$705 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$210 \$706 \$147 \$177 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$211 \$180 \$304 \$706 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$212 \$179 \$303 \$180 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$213 b5_r7_b_not \$303 \$84 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$214 \$707 \$304 b5_r7_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$215 \$180 \$147 \$707 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$216 \$708 \$147 \$84 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$217 b5_r7_b \$304 \$708 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$218 \$180 \$303 b5_r7_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$219 \$184 b6|b6_q0|b6_q1|b6_q2|b6_q3|b6_q4|b6_q5|b6_q6|b6_q7 b6_c7_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$220 \$709
+ b6_not|b6_q0_not|b6_q1_not|b6_q2_not|b6_q3_not|b6_q4_not|b6_q5_not|b6_q6_not|b6_q7_not
+ \$184 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$221 b6_c7
+ a7_not|b0_p7_not|b1_p7_not|b2_p7_not|b4_p7_not|b5_p7_not|b6_p7_not|b7_p7_not
+ \$709 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$222 \$710
+ a7_not|b0_p7_not|b1_p7_not|b2_p7_not|b4_p7_not|b5_p7_not|b6_p7_not|b7_p7_not
+ b6_c7_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$223 \$186
+ b6_not|b6_q0_not|b6_q1_not|b6_q2_not|b6_q3_not|b6_q4_not|b6_q5_not|b6_q6_not|b6_q7_not
+ \$710 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$224 b6_c7 b6|b6_q0|b6_q1|b6_q2|b6_q3|b6_q4|b6_q5|b6_q6|b6_q7 \$186 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$225 \$86 \$311 \$184 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$226 \$711 \$312 \$86 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$227 \$186 \$148 \$711 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$228 \$712 \$148 \$184 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$229 \$187 \$312 \$712 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$230 \$186 \$311 \$187 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$231 b6_r7_b_not \$311 \$86 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$232 \$713 \$312 b6_r7_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$233 \$187 \$148 \$713 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$234 \$714 \$148 \$86 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$235 b6_r7_b \$312 \$714 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$236 \$187 \$311 b6_r7_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$237 \$191 b1_q3|b7|b7_q0|b7_q1|b7_q2|b7_q4|b7_q5|b7_q6|b7_q7 b6_c7_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$238 \$715
+ b7_not|b7_q0_not|b7_q1_not|b7_q2_not|b7_q3_not|b7_q4_not|b7_q5_not|b7_q6_not|b7_q7_not
+ \$191 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$239 b6_c7
+ a7_not|b0_p7_not|b1_p7_not|b2_p7_not|b4_p7_not|b5_p7_not|b6_p7_not|b7_p7_not
+ \$715 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$240 \$716
+ a7_not|b0_p7_not|b1_p7_not|b2_p7_not|b4_p7_not|b5_p7_not|b6_p7_not|b7_p7_not
+ b6_c7_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$241 \$193
+ b7_not|b7_q0_not|b7_q1_not|b7_q2_not|b7_q3_not|b7_q4_not|b7_q5_not|b7_q6_not|b7_q7_not
+ \$716 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$242 b6_c7 b1_q3|b7|b7_q0|b7_q1|b7_q2|b7_q4|b7_q5|b7_q6|b7_q7 \$193 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$243 \$88 \$319 \$191 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$244 \$717 \$320 \$88 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$245 \$193 \$149 \$717 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$246 \$718 \$149 \$191 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$247 \$194 \$320 \$718 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$248 \$193 \$319 \$194 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$249 \$195 \$319 \$88 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$250 \$719 \$320 \$195 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$251 \$194 \$149 \$719 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$252 \$720 \$149 \$88 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$253 \$196 \$320 \$720 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$254 \$194 \$319 \$196 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$255 \$1397 b1|b1_q0|b1_q1|b1_q2|b1_q3|b1_q4|b1_q5|b1_q6|b1_q7 b1_c6_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$256 \$220 a7|b0_p7|b1_p7|b2_p7|b3_p7|b4_p7|b5_p7|b6_p7|b7_p7 b1_c7_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$257 \$1637
+ b1_not|b1_q0_not|b1_q1_not|b1_q2_not|b1_q3_not|b1_q4_not|b1_q5_not|b1_q6_not|b1_q7_not
+ \$1397 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$258 b1_c6
+ a6_not|b0_p6_not|b1_p6_not|b3_p6_not|b4_p6_not|b5_p6_not|b6_p6_not|b7_p6_not
+ \$1637 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$259 \$1638
+ a6_not|b0_p6_not|b1_p6_not|b3_p6_not|b4_p6_not|b5_p6_not|b6_p6_not|b7_p6_not
+ b1_c6_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$260 \$1107
+ b1_not|b1_q0_not|b1_q1_not|b1_q2_not|b1_q3_not|b1_q4_not|b1_q5_not|b1_q6_not|b1_q7_not
+ \$1638 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$261 b1_c6 b1|b1_q0|b1_q1|b1_q2|b1_q3|b1_q4|b1_q5|b1_q6|b1_q7 \$1107 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$262 b1_c7 a7|b0_p7|b1_p7|b2_p7|b3_p7|b4_p7|b5_p7|b6_p7|b7_p7 \$151 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$263 \$1252 \$1110 \$1397 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$264 \$1107 \$1112 \$1252 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$265 \$1253 \$1110 \$1107 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$266 \$1397 \$1112 \$1253 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$267 \$1254 \$1110 \$1402 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$268 \$1403 \$1112 \$1254 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$269 \$725 \$1110 \$1403 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$270 \$1402 \$1112 \$725 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$271 \$76 \$273 x0_a7_f_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$272 x0_a7_f \$273 \$152 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$273 x0_a7_b_not \$273 \$76 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$274 b0_r7_b_not \$1252 \$275 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$275 \$1643 \$1253 b0_r7_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$276 \$274 \$725 \$1643 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$277 \$1644 \$725 \$275 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$278 b0_r7_b \$1253 \$1644 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$279 \$152 \$273 x0_a7_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$280 \$274 \$1252 b0_r7_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$281 \$1190 b0_r7_b_not \$725 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$282 \$1254 b0_r7_b \$1190 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$283 \$1191 b0_r7_b_not \$1254 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$284 \$725 b0_r7_b \$1191 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$285 \$1192 \$1191 \$1253 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$286 \$1252 \$1190 \$1192 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$287 \$1193 \$1191 \$1252 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$288 \$1253 \$1190 \$1193 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$289 \$156 a7|b0_p7|b1_p7|b2_p7|b3_p7|b4_p7|b5_p7|b6_p7|b7_p7 b2_c7_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$290 b2_c7 a7|b0_p7|b1_p7|b2_p7|b3_p7|b4_p7|b5_p7|b6_p7|b7_p7 \$158 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$291 \$1257 \$1117 \$277 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$292 \$276 \$1119 \$1257 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$293 \$1258 \$1117 \$276 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$294 \$277 \$1119 \$1258 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$295 \$1259 \$1117 \$1411 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$296 \$1412 \$1119 \$1259 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$297 \$727 \$1117 \$1412 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$298 \$1411 \$1119 \$727 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$299 \$78 \$281 \$156 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$300 \$158 \$281 \$159 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$301 b2_r6_b_not \$1257 \$283 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$302 b2_r7_b_not \$281 \$78 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$303 \$1649 \$1258 b2_r6_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$304 \$282 \$727 \$1649 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$305 \$1650 \$727 \$283 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$306 b2_r6_b \$1258 \$1650 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$307 \$159 \$281 b2_r7_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$308 \$282 \$1257 b2_r6_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$309 \$1194 b2_r6_b_not \$727 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$310 \$1259 b2_r6_b \$1194 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$311 \$1195 b2_r6_b_not \$1259 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$312 \$727 b2_r6_b \$1195 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$313 \$1196 \$1195 \$1258 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$314 \$1257 \$1194 \$1196 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$315 \$1197 \$1195 \$1257 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$316 \$1258 \$1194 \$1197 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$317 \$163 a7|b0_p7|b1_p7|b2_p7|b3_p7|b4_p7|b5_p7|b6_p7|b7_p7 b3_c7_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$318 \$1123
+ b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b3|b3_q0|b3_q1|b3_q2|b3_q3|b3_q4|b3_q5|b3_q6|b3_q7
+ b3_c6_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$319 \$1651
+ b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b3_not|b3_q0_not|b3_q1_not|b3_q2_not|b3_q3_not|b3_q4_not|b3_q5_not|b3_q6_not|b3_q7_not
+ \$1123 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$320 b3_c6
+ a6_not|b0_p6_not|b1_p6_not|b3_p6_not|b4_p6_not|b5_p6_not|b6_p6_not|b7_p6_not
+ \$1651 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$321 \$1652
+ a6_not|b0_p6_not|b1_p6_not|b3_p6_not|b4_p6_not|b5_p6_not|b6_p6_not|b7_p6_not
+ b3_c6_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$322 \$1125
+ b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b3_not|b3_q0_not|b3_q1_not|b3_q2_not|b3_q3_not|b3_q4_not|b3_q5_not|b3_q6_not|b3_q7_not
+ \$1652 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$323 b3_c7 a7|b0_p7|b1_p7|b2_p7|b3_p7|b4_p7|b5_p7|b6_p7|b7_p7 \$165 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$324 b3_c6
+ b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b3|b3_q0|b3_q1|b3_q2|b3_q3|b3_q4|b3_q5|b3_q6|b3_q7
+ \$1125 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$325 \$1198 \$1123 \$285 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$326 \$284 \$1125 \$1198 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$327 \$1199 \$1123 \$284 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$328 \$285 \$1125 \$1199 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$329 \$1200 \$1123 \$1420 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$330 \$1421 \$1125 \$1200 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$331 \$729 \$1123 \$1421 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$332 \$1420 \$1125 \$729 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$333 \$80 \$288 \$163 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$334 \$223 \$1198 \$1123 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$335 \$1653 \$1199 \$223 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$336 \$1125 \$729 \$1653 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$337 \$1654 \$729 \$1123 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$338 \$451 \$1199 \$1654 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$339 \$165 \$288 \$166 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$340 \$1125 \$1198 \$451 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$341 b3_r7_b_not \$288 \$80 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$342 b3_r6_b_not \$1198 \$291 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$343 \$1655 \$1199 b3_r6_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$344 \$290 \$729 \$1655 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$345 \$1656 \$729 \$291 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$346 b3_r6_b \$1199 \$1656 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$347 \$166 \$288 b3_r7_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$348 \$290 \$1198 b3_r6_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$349 \$1201 b3_r6_b_not \$729 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$350 \$1200 b3_r6_b \$1201 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$351 \$1202 b3_r6_b_not \$1200 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$352 \$729 b3_r6_b \$1202 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$353 \$1203 \$1202 \$1199 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$354 \$1198 \$1201 \$1203 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$355 \$1204 \$1202 \$1198 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$356 \$1199 \$1201 \$1204 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$357 \$170 a7|b0_p7|b1_p7|b2_p7|b3_p7|b4_p7|b5_p7|b6_p7|b7_p7 b4_c7_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$358 \$170 b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b4|b4_q7 b4_c7_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$359 \$730
+ b2_q0_not|b2_q1_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b4_not|b4_q7_not
+ \$170 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$360 b4_c7
+ a7_not|b0_p7_not|b1_p7_not|b2_p7_not|b4_p7_not|b5_p7_not|b6_p7_not|b7_p7_not
+ \$730 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$361 \$731
+ a7_not|b0_p7_not|b1_p7_not|b2_p7_not|b4_p7_not|b5_p7_not|b6_p7_not|b7_p7_not
+ b4_c7_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$362 \$172
+ b2_q0_not|b2_q1_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b4_not|b4_q7_not
+ \$731 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$363 b4_c7 b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b4|b4_q7 \$172 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$364 b4_c7 a7|b0_p7|b1_p7|b2_p7|b3_p7|b4_p7|b5_p7|b6_p7|b7_p7 \$172 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$365 \$1264 \$1129 \$293 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$366 \$292 \$1131 \$1264 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$367 \$1265 \$1129 \$292 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$368 \$293 \$1131 \$1265 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$369 \$1266 \$1129 \$1429 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$370 \$1430 \$1131 \$1266 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$371 \$733 \$1129 \$1430 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$372 \$1429 \$1131 \$733 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$373 \$82 \$297 \$170 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$374 \$172 \$297 \$173 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$375 b4_r6_b_not \$1264 \$299 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$376 b4_r7_b_not \$297 \$82 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$377 \$1661 \$1265 b4_r6_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$378 \$298 \$733 \$1661 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$379 \$1662 \$733 \$299 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$380 b4_r6_b \$1265 \$1662 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$381 \$298 \$1264 b4_r6_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$382 \$173 \$297 b4_r7_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$383 \$1205 b4_r6_b_not \$733 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$384 \$1266 b4_r6_b \$1205 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$385 \$1206 b4_r6_b_not \$1266 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$386 \$733 b4_r6_b \$1206 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$387 \$1207 \$1206 \$1265 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$388 \$1264 \$1205 \$1207 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$389 \$1208 \$1206 \$1264 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$390 \$1265 \$1205 \$1208 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$391 \$177 a7|b0_p7|b1_p7|b2_p7|b3_p7|b4_p7|b5_p7|b6_p7|b7_p7 b5_c7_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$392 \$177 b5|b5_q0|b5_q1|b5_q2|b5_q3|b5_q4|b5_q5|b5_q6|b5_q7 b5_c7_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$393 \$734
+ b5_not|b5_q0_not|b5_q1_not|b5_q2_not|b5_q3_not|b5_q4_not|b5_q5_not|b5_q6_not|b5_q7_not
+ \$177 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$394 b5_c7
+ a7_not|b0_p7_not|b1_p7_not|b2_p7_not|b4_p7_not|b5_p7_not|b6_p7_not|b7_p7_not
+ \$734 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$395 \$735
+ a7_not|b0_p7_not|b1_p7_not|b2_p7_not|b4_p7_not|b5_p7_not|b6_p7_not|b7_p7_not
+ b5_c7_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$396 \$179
+ b5_not|b5_q0_not|b5_q1_not|b5_q2_not|b5_q3_not|b5_q4_not|b5_q5_not|b5_q6_not|b5_q7_not
+ \$735 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$397 b5_c7 b5|b5_q0|b5_q1|b5_q2|b5_q3|b5_q4|b5_q5|b5_q6|b5_q7 \$179 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$398 b5_c7 a7|b0_p7|b1_p7|b2_p7|b3_p7|b4_p7|b5_p7|b6_p7|b7_p7 \$179 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$399 \$1269 \$1135 \$301 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$400 \$300 \$1137 \$1269 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$401 \$1270 \$1135 \$300 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$402 \$301 \$1137 \$1270 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$403 \$1271 \$1135 \$1438 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$404 \$1439 \$1137 \$1271 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$405 \$737 \$1135 \$1439 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$406 \$1438 \$1137 \$737 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$407 \$84 \$305 \$177 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$408 \$179 \$305 \$180 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$409 b5_r6_b_not \$1269 \$307 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$410 b5_r7_b_not \$305 \$84 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$411 \$1667 \$1270 b5_r6_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$412 \$306 \$737 \$1667 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$413 \$1668 \$737 \$307 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$414 b5_r6_b \$1270 \$1668 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$415 \$306 \$1269 b5_r6_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$416 \$180 \$305 b5_r7_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$417 \$1209 b5_r6_b_not \$737 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$418 \$1271 b5_r6_b \$1209 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$419 \$1210 b5_r6_b_not \$1271 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$420 \$737 b5_r6_b \$1210 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$421 \$1211 \$1210 \$1270 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$422 \$1269 \$1209 \$1211 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$423 \$1212 \$1210 \$1269 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$424 \$1270 \$1209 \$1212 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$425 \$184 a7|b0_p7|b1_p7|b2_p7|b3_p7|b4_p7|b5_p7|b6_p7|b7_p7 b6_c7_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$426 b6_c7 a7|b0_p7|b1_p7|b2_p7|b3_p7|b4_p7|b5_p7|b6_p7|b7_p7 \$186 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$427 \$1274 \$1141 \$309 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$428 \$308 \$1143 \$1274 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$429 \$1275 \$1141 \$308 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$430 \$309 \$1143 \$1275 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$431 \$1276 \$1141 \$1447 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$432 \$1448 \$1143 \$1276 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$433 \$739 \$1141 \$1448 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$434 \$1447 \$1143 \$739 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$435 \$86 \$313 \$184 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$436 \$186 \$313 \$187 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$437 b6_r7_b_not \$313 \$86 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$438 b6_r6_b_not \$1274 \$315 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$439 \$1673 \$1275 b6_r6_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$440 \$314 \$739 \$1673 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$441 \$1674 \$739 \$315 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$442 b6_r6_b \$1275 \$1674 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$443 \$314 \$1274 b6_r6_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$444 \$187 \$313 b6_r7_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$445 \$1213 b6_r6_b_not \$739 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$446 \$1276 b6_r6_b \$1213 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$447 \$1214 b6_r6_b_not \$1276 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$448 \$739 b6_r6_b \$1214 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$449 \$1215 \$1214 \$1275 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$450 \$1274 \$1213 \$1215 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$451 \$1216 \$1214 \$1274 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$452 \$1275 \$1213 \$1216 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$453 \$191 a7|b0_p7|b1_p7|b2_p7|b3_p7|b4_p7|b5_p7|b6_p7|b7_p7 b6_c7_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$454 b6_c7 a7|b0_p7|b1_p7|b2_p7|b3_p7|b4_p7|b5_p7|b6_p7|b7_p7 \$193 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$455 \$1279 \$1147 \$317 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$456 \$316 \$1149 \$1279 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$457 \$1280 \$1147 \$316 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$458 \$317 \$1149 \$1280 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$459 \$1281 \$1147 \$1456 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$460 \$1457 \$1149 \$1281 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$461 \$741 \$1147 \$1457 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$462 \$1456 \$1149 \$741 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$463 \$88 \$321 \$191 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$464 \$193 \$321 \$194 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$465 \$195 \$321 \$88 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$466 \$1150 \$1279 \$323 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$467 \$1679 \$1280 \$1150 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$468 \$322 \$741 \$1679 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$469 \$1680 \$741 \$323 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$470 \$1151 \$1280 \$1680 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$471 \$194 \$321 \$196 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$472 \$322 \$1279 \$1151 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$473 \$1217 \$1150 \$741 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$474 \$1281 \$1151 \$1217 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$475 \$1218 \$1150 \$1281 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$476 \$741 \$1151 \$1218 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$477 p13 \$1218 \$1280 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$478 \$1279 \$1217 p13 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$479 p13_not \$1218 \$1279 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$480 \$1280 \$1217 p13_not vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$481 \$1397 a6|b0_p6|b1_p6|b3_p6|b4_p6|b5_p6|b6_p6|b7_p6 b1_c6_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$482 b1_c6 a6|b0_p6|b1_p6|b3_p6|b4_p6|b5_p6|b6_p6|b7_p6 \$1107 vdd pfet_03v3
+ L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$483 \$1110 a7|b0_p7|b1_p7|b2_p7|b3_p7|b4_p7|b5_p7|b6_p7|b7_p7 b0_c7_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$484 \$1110 b0|b0_q0|b0_q1|b0_q2|b0_q3|b0_q4|b0_q5|b0_q6|b0_q7 b0_c7_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$485 \$1639
+ b0_not|b0_q0_not|b0_q1_not|b0_q3_not|b0_q4_not|b0_q5_not|b0_q6_not|b0_q7_not|b1_q2_not
+ \$1110 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$486 b0_c7
+ a7_not|b0_p7_not|b1_p7_not|b2_p7_not|b4_p7_not|b5_p7_not|b6_p7_not|b7_p7_not
+ \$1639 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$487 \$1640
+ a7_not|b0_p7_not|b1_p7_not|b2_p7_not|b4_p7_not|b5_p7_not|b6_p7_not|b7_p7_not
+ b0_c7_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$488 \$1112
+ b0_not|b0_q0_not|b0_q1_not|b0_q3_not|b0_q4_not|b0_q5_not|b0_q6_not|b0_q7_not|b1_q2_not
+ \$1640 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$489 b0_c7 a7|b0_p7|b1_p7|b2_p7|b3_p7|b4_p7|b5_p7|b6_p7|b7_p7 \$1112 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$490 b0_c7 b0|b0_q0|b0_q1|b0_q2|b0_q3|b0_q4|b0_q5|b0_q6|b0_q7 \$1112 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$491 \$2208 \$2085 \$2358 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$492 \$2358 \$2086 \$2210 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$493 \$2209 \$2085 \$2360 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$494 \$2360 \$2086 \$2068 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$495 \$221 \$1254 \$1110 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$496 \$221 \$1252 \$1110 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$497 \$1641 \$1253 \$221 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$498 \$1112 \$725 \$1641 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$499 \$1642 \$725 \$1110 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$500 \$608 \$1253 \$1642 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$501 \$1112 \$1252 \$608 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$502 \$1112 \$1254 \$608 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$503 b0_r7_b_not \$1254 \$275 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$504 \$274 \$1254 b0_r7_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$505 \$1117 a6|b0_p6|b1_p6|b3_p6|b4_p6|b5_p6|b6_p6|b7_p6 b2_c6_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$506 \$1117 b2|b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7 b2_c6_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$507 \$1645
+ b2_not|b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not
+ \$1117 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$508 b2_c6
+ a6_not|b0_p6_not|b1_p6_not|b3_p6_not|b4_p6_not|b5_p6_not|b6_p6_not|b7_p6_not
+ \$1645 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$509 \$1646
+ a6_not|b0_p6_not|b1_p6_not|b3_p6_not|b4_p6_not|b5_p6_not|b6_p6_not|b7_p6_not
+ b2_c6_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$510 \$1119
+ b2_not|b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not
+ \$1646 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$511 b2_c6 a6|b0_p6|b1_p6|b3_p6|b4_p6|b5_p6|b6_p6|b7_p6 \$1119 vdd pfet_03v3
+ L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$512 b2_c6 b2|b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7 \$1119 vdd pfet_03v3
+ L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$513 \$2215 \$2090 \$1193 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$514 \$1193 \$2091 \$2217 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$515 \$2216 \$2090 \$2368 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$516 \$2368 \$2091 \$2070 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$517 \$222 \$1257 \$1117 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$518 \$222 \$1259 \$1117 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$519 \$1647 \$1258 \$222 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$520 \$1119 \$727 \$1647 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$521 \$1648 \$727 \$1117 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$522 \$613 \$1258 \$1648 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$523 \$1119 \$1259 \$613 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$524 \$1119 \$1257 \$613 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$525 b2_r6_b_not \$1259 \$283 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$526 \$282 \$1259 b2_r6_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$527 \$1123 a6|b0_p6|b1_p6|b3_p6|b4_p6|b5_p6|b6_p6|b7_p6 b3_c6_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$528 b3_c6 a6|b0_p6|b1_p6|b3_p6|b4_p6|b5_p6|b6_p6|b7_p6 \$1125 vdd pfet_03v3
+ L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$529 \$2162 \$2095 \$1197 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$530 \$1196 \$2096 \$2162 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$531 \$2163 \$2095 \$1196 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$532 \$1197 \$2096 \$2163 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$533 \$2164 \$2095 \$2375 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$534 \$2376 \$2096 \$2164 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$535 \$2072 \$2095 \$2376 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$536 \$2375 \$2096 \$2072 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$537 \$223 \$1200 \$1123 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$538 \$1125 \$1200 \$451 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$539 b3_r6_b_not \$1200 \$291 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$540 \$290 \$1200 b3_r6_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$541 \$2165 b3_r5_b_not \$2072 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$542 \$2164 b3_r5_b \$2165 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$543 \$2072 b3_r5_b \$2166 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$544 \$2167 \$2166 \$2163 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$545 \$2162 \$2165 \$2167 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$546 \$2163 \$2165 \$2168 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$547 \$1129 b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b4|b4_q7 b4_c6_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$548 \$1129 a6|b0_p6|b1_p6|b3_p6|b4_p6|b5_p6|b6_p6|b7_p6 b4_c6_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$549 \$1657
+ b2_q0_not|b2_q1_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b4_not|b4_q7_not
+ \$1129 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$550 b4_c6
+ a6_not|b0_p6_not|b1_p6_not|b3_p6_not|b4_p6_not|b5_p6_not|b6_p6_not|b7_p6_not
+ \$1657 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$551 \$1658
+ a6_not|b0_p6_not|b1_p6_not|b3_p6_not|b4_p6_not|b5_p6_not|b6_p6_not|b7_p6_not
+ b4_c6_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$552 \$1131
+ b2_q0_not|b2_q1_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b4_not|b4_q7_not
+ \$1658 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$553 b4_c6 b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b4|b4_q7 \$1131 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$554 b4_c6 a6|b0_p6|b1_p6|b3_p6|b4_p6|b5_p6|b6_p6|b7_p6 \$1131 vdd pfet_03v3
+ L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$555 \$2169 \$2100 \$1204 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$556 \$1203 \$2101 \$2169 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$557 \$1204 \$2101 \$2224 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$558 \$2170 \$2100 \$2383 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$559 \$2384 \$2101 \$2170 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$560 \$2383 \$2101 \$2074 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$561 \$224 \$1266 \$1129 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$562 \$224 \$1264 \$1129 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$563 \$1659 \$1265 \$224 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$564 \$1131 \$733 \$1659 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$565 \$1660 \$733 \$1129 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$566 \$622 \$1265 \$1660 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$567 \$1131 \$1266 \$622 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$568 \$1131 \$1264 \$622 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$569 b4_r6_b_not \$1266 \$299 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$570 \$298 \$1266 b4_r6_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$571 \$2225 b4_r5_b_not \$2074 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$572 \$2074 b4_r5_b \$2226 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$573 \$2227 \$2226 \$2224 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$574 \$2224 \$2225 \$2228 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$575 \$1135 b5|b5_q0|b5_q1|b5_q2|b5_q3|b5_q4|b5_q5|b5_q6|b5_q7 b5_c6_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$576 \$1135 a6|b0_p6|b1_p6|b3_p6|b4_p6|b5_p6|b6_p6|b7_p6 b5_c6_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$577 \$1663
+ b5_not|b5_q0_not|b5_q1_not|b5_q2_not|b5_q3_not|b5_q4_not|b5_q5_not|b5_q6_not|b5_q7_not
+ \$1135 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$578 b5_c6
+ a6_not|b0_p6_not|b1_p6_not|b3_p6_not|b4_p6_not|b5_p6_not|b6_p6_not|b7_p6_not
+ \$1663 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$579 \$1664
+ a6_not|b0_p6_not|b1_p6_not|b3_p6_not|b4_p6_not|b5_p6_not|b6_p6_not|b7_p6_not
+ b5_c6_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$580 \$1137
+ b5_not|b5_q0_not|b5_q1_not|b5_q2_not|b5_q3_not|b5_q4_not|b5_q5_not|b5_q6_not|b5_q7_not
+ \$1664 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$581 b5_c6 b5|b5_q0|b5_q1|b5_q2|b5_q3|b5_q4|b5_q5|b5_q6|b5_q7 \$1137 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$582 b5_c6 a6|b0_p6|b1_p6|b3_p6|b4_p6|b5_p6|b6_p6|b7_p6 \$1137 vdd pfet_03v3
+ L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$583 \$2171 \$2106 \$1208 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$584 \$1207 \$2107 \$2171 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$585 \$1208 \$2107 \$2229 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$586 \$2172 \$2106 \$2391 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$587 \$2392 \$2107 \$2172 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$588 \$2391 \$2107 \$2076 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$589 \$225 \$1271 \$1135 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$590 \$225 \$1269 \$1135 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$591 \$1665 \$1270 \$225 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$592 \$1137 \$737 \$1665 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$593 \$1666 \$737 \$1135 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$594 \$627 \$1270 \$1666 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$595 \$1137 \$1269 \$627 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$596 \$1137 \$1271 \$627 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$597 b5_r6_b_not \$1271 \$307 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$598 \$306 \$1271 b5_r6_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$599 \$2230 b5_r5_b_not \$2076 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$600 \$2076 b5_r5_b \$2231 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$601 \$2232 \$2231 \$2229 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$602 \$2229 \$2230 \$2233 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$603 \$1141 a6|b0_p6|b1_p6|b3_p6|b4_p6|b5_p6|b6_p6|b7_p6 b6_c6_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$604 \$1141 b6|b6_q0|b6_q1|b6_q2|b6_q3|b6_q4|b6_q5|b6_q6|b6_q7 b6_c6_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$605 \$1669
+ b6_not|b6_q0_not|b6_q1_not|b6_q2_not|b6_q3_not|b6_q4_not|b6_q5_not|b6_q6_not|b6_q7_not
+ \$1141 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$606 b6_c6
+ a6_not|b0_p6_not|b1_p6_not|b3_p6_not|b4_p6_not|b5_p6_not|b6_p6_not|b7_p6_not
+ \$1669 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$607 \$1670
+ a6_not|b0_p6_not|b1_p6_not|b3_p6_not|b4_p6_not|b5_p6_not|b6_p6_not|b7_p6_not
+ b6_c6_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$608 \$1143
+ b6_not|b6_q0_not|b6_q1_not|b6_q2_not|b6_q3_not|b6_q4_not|b6_q5_not|b6_q6_not|b6_q7_not
+ \$1670 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$609 b6_c6 b6|b6_q0|b6_q1|b6_q2|b6_q3|b6_q4|b6_q5|b6_q6|b6_q7 \$1143 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$610 b6_c6 a6|b0_p6|b1_p6|b3_p6|b4_p6|b5_p6|b6_p6|b7_p6 \$1143 vdd pfet_03v3
+ L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$611 \$2173 \$2111 \$1212 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$612 \$1211 \$2112 \$2173 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$613 \$1212 \$2112 \$2236 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$614 \$2174 \$2111 \$2398 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$615 \$2399 \$2112 \$2174 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$616 \$2398 \$2112 \$2078 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$617 \$226 \$1274 \$1141 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$618 \$226 \$1276 \$1141 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$619 \$1671 \$1275 \$226 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$620 \$1143 \$739 \$1671 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$621 \$1672 \$739 \$1141 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$622 \$632 \$1275 \$1672 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$623 \$1143 \$1276 \$632 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$624 \$1143 \$1274 \$632 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$625 b6_r6_b_not \$1276 \$315 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$626 \$314 \$1276 b6_r6_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$627 \$2237 b6_r5_b_not \$2078 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$628 \$2078 b6_r5_b \$2238 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$629 \$2239 \$2238 \$2236 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$630 \$2236 \$2237 \$2240 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$631 \$1147 b1_q3|b7|b7_q0|b7_q1|b7_q2|b7_q4|b7_q5|b7_q6|b7_q7 b6_c6_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$632 \$1147 a6|b0_p6|b1_p6|b3_p6|b4_p6|b5_p6|b6_p6|b7_p6 b6_c6_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$633 \$1675
+ b7_not|b7_q0_not|b7_q1_not|b7_q2_not|b7_q3_not|b7_q4_not|b7_q5_not|b7_q6_not|b7_q7_not
+ \$1147 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$634 b6_c6
+ a6_not|b0_p6_not|b1_p6_not|b3_p6_not|b4_p6_not|b5_p6_not|b6_p6_not|b7_p6_not
+ \$1675 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$635 \$1676
+ a6_not|b0_p6_not|b1_p6_not|b3_p6_not|b4_p6_not|b5_p6_not|b6_p6_not|b7_p6_not
+ b6_c6_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$636 \$1149
+ b7_not|b7_q0_not|b7_q1_not|b7_q2_not|b7_q3_not|b7_q4_not|b7_q5_not|b7_q6_not|b7_q7_not
+ \$1676 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$637 b6_c6 b1_q3|b7|b7_q0|b7_q1|b7_q2|b7_q4|b7_q5|b7_q6|b7_q7 \$1149 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$638 b6_c6 a6|b0_p6|b1_p6|b3_p6|b4_p6|b5_p6|b6_p6|b7_p6 \$1149 vdd pfet_03v3
+ L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$639 \$2175 \$2116 \$1216 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$640 \$1215 \$2117 \$2175 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$641 \$1216 \$2117 \$2241 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$642 \$2176 \$2116 \$2406 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$643 \$2407 \$2117 \$2176 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$644 \$2406 \$2117 \$2080 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$645 \$227 \$1279 \$1147 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$646 \$227 \$1281 \$1147 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$647 \$1677 \$1280 \$227 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$648 \$1149 \$741 \$1677 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$649 \$1678 \$741 \$1147 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$650 \$637 \$1280 \$1678 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$651 \$1149 \$1281 \$637 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$652 \$1149 \$1279 \$637 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$653 \$1150 \$1281 \$323 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$654 \$322 \$1281 \$1151 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$655 \$2242 \$2118 \$2080 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$656 \$2080 \$2119 \$2243 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$657 p12 \$2243 \$2241 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$658 \$2241 \$2242 p12_not vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$659 \$2358 b1|b1_q0|b1_q1|b1_q2|b1_q3|b1_q4|b1_q5|b1_q6|b1_q7 b1_c5_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$660 \$2603
+ b1_not|b1_q0_not|b1_q1_not|b1_q2_not|b1_q3_not|b1_q4_not|b1_q5_not|b1_q6_not|b1_q7_not
+ \$2358 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$661 b1_c5
+ a5_not|b0_p5_not|b1_p5_not|b2_p5_not|b3_p5_not|b5_p5_not|b6_p5_not|b7_p5_not
+ \$2603 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$662 \$2604
+ a5_not|b0_p5_not|b1_p5_not|b2_p5_not|b3_p5_not|b5_p5_not|b6_p5_not|b7_p5_not
+ b1_c5_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$663 \$2083
+ b1_not|b1_q0_not|b1_q1_not|b1_q2_not|b1_q3_not|b1_q4_not|b1_q5_not|b1_q6_not|b1_q7_not
+ \$2604 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$664 b1_c5 b1|b1_q0|b1_q1|b1_q2|b1_q3|b1_q4|b1_q5|b1_q6|b1_q7 \$2083 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$665 \$2083 \$2086 \$2208 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$666 \$2210 \$2085 \$2083 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$667 \$2361 \$2086 \$2209 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$668 \$2068 \$2085 \$2361 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$669 \$2211 b0_r6_b_not \$2068 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$670 \$2209 b0_r6_b \$2211 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$671 \$2212 b0_r6_b_not \$2209 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$672 \$2068 b0_r6_b \$2212 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$673 \$2213 \$2212 \$2210 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$674 \$2208 \$2211 \$2213 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$675 \$2214 \$2212 \$2208 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$676 \$2210 \$2211 \$2214 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$677 \$1192 \$2091 \$2215 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$678 \$2217 \$2090 \$1192 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$679 \$2369 \$2091 \$2216 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$680 \$2070 \$2090 \$2369 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$681 \$2218 b2_r5_b_not \$2070 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$682 \$2216 b2_r5_b \$2218 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$683 \$2219 b2_r5_b_not \$2216 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$684 \$2070 b2_r5_b \$2219 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$685 \$2220 \$2219 \$2217 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$686 \$2215 \$2218 \$2220 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$687 \$2221 \$2219 \$2215 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$688 \$2217 \$2218 \$2221 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$689 \$2095
+ b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b3|b3_q0|b3_q1|b3_q2|b3_q3|b3_q4|b3_q5|b3_q6|b3_q7
+ b2_c5_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$690 \$2617
+ b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b3_not|b3_q0_not|b3_q1_not|b3_q2_not|b3_q3_not|b3_q4_not|b3_q5_not|b3_q6_not|b3_q7_not
+ \$2095 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$691 b3_c5
+ a5_not|b0_p5_not|b1_p5_not|b2_p5_not|b3_p5_not|b5_p5_not|b6_p5_not|b7_p5_not
+ \$2617 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$692 \$2618
+ a5_not|b0_p5_not|b1_p5_not|b2_p5_not|b3_p5_not|b5_p5_not|b6_p5_not|b7_p5_not
+ b2_c5_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$693 \$2096
+ b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b3_not|b3_q0_not|b3_q1_not|b3_q2_not|b3_q3_not|b3_q4_not|b3_q5_not|b3_q6_not|b3_q7_not
+ \$2618 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$694 b3_c5
+ b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b3|b3_q0|b3_q1|b3_q2|b3_q3|b3_q4|b3_q5|b3_q6|b3_q7
+ \$2096 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$695 \$2166 b3_r5_b_not \$2164 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$696 \$2168 \$2166 \$2162 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$697 \$2224 \$2100 \$1203 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$698 \$2074 \$2100 \$2384 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$699 \$2170 b4_r5_b \$2225 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$700 \$2226 b4_r5_b_not \$2170 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$701 \$2169 \$2225 \$2227 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$702 \$2228 \$2226 \$2169 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$703 \$2229 \$2106 \$1207 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$704 \$2076 \$2106 \$2392 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$705 \$2172 b5_r5_b \$2230 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$706 \$2231 b5_r5_b_not \$2172 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$707 \$2171 \$2230 \$2232 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$708 \$2233 \$2231 \$2171 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$709 \$2236 \$2111 \$1211 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$710 \$2078 \$2111 \$2399 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$711 \$2174 b6_r5_b \$2237 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$712 \$2238 b6_r5_b_not \$2174 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$713 \$2173 \$2237 \$2239 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$714 \$2240 \$2238 \$2173 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$715 \$2241 \$2116 \$1215 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$716 \$2080 \$2116 \$2407 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$717 \$2176 \$2119 \$2242 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$718 \$2243 \$2118 \$2176 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$719 \$2175 \$2242 p12 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$720 p12_not \$2243 \$2175 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$721 \$2358 a5|b0_p5|b1_p5|b3_p5|b4_p5|b5_p5|b6_p5|b7_p5 b1_c5_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$722 \$2085 a6|b0_p6|b1_p6|b3_p6|b4_p6|b5_p6|b6_p6|b7_p6 b0_c6_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$723 \$2085 b0|b0_q0|b0_q1|b0_q2|b0_q3|b0_q4|b0_q5|b0_q6|b0_q7 b0_c6_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$724 \$2605
+ b0_not|b0_q0_not|b0_q1_not|b0_q3_not|b0_q4_not|b0_q5_not|b0_q6_not|b0_q7_not|b1_q2_not
+ \$2085 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$725 b0_c6
+ a6_not|b0_p6_not|b1_p6_not|b3_p6_not|b4_p6_not|b5_p6_not|b6_p6_not|b7_p6_not
+ \$2605 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$726 \$2606
+ a6_not|b0_p6_not|b1_p6_not|b3_p6_not|b4_p6_not|b5_p6_not|b6_p6_not|b7_p6_not
+ b0_c6_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$727 \$2086
+ b0_not|b0_q0_not|b0_q1_not|b0_q3_not|b0_q4_not|b0_q5_not|b0_q6_not|b0_q7_not|b1_q2_not
+ \$2606 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$728 b0_c6 b0|b0_q0|b0_q1|b0_q2|b0_q3|b0_q4|b0_q5|b0_q6|b0_q7 \$2086 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$729 \$1402 \$2208 \$2085 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$730 \$2607 \$2210 \$1402 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$731 \$2086 \$2068 \$2607 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$732 \$2608 \$2068 \$2085 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$733 \$1403 \$2210 \$2608 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$734 \$2086 \$2208 \$1403 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$735 b0_r6_b_not \$2208 \$1191 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$736 \$2609 \$2210 b0_r6_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$737 \$1190 \$2068 \$2609 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$738 \$2610 \$2068 \$1191 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$739 b0_r6_b \$2210 \$2610 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$740 \$1190 \$2208 b0_r6_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$741 \$2090 b2|b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7 b2_c5_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$742 \$2611
+ b2_not|b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not
+ \$2090 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$743 b2_c5
+ a5_not|b0_p5_not|b1_p5_not|b2_p5_not|b3_p5_not|b5_p5_not|b6_p5_not|b7_p5_not
+ \$2611 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$744 \$2612
+ a5_not|b0_p5_not|b1_p5_not|b2_p5_not|b3_p5_not|b5_p5_not|b6_p5_not|b7_p5_not
+ b2_c5_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$745 \$2091
+ b2_not|b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not
+ \$2612 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$746 b2_c5 b2|b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7 \$2091 vdd pfet_03v3
+ L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$747 \$1411 \$2215 \$2090 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$748 \$2613 \$2217 \$1411 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$749 \$2091 \$2070 \$2613 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$750 \$2614 \$2070 \$2090 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$751 \$1412 \$2217 \$2614 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$752 \$2091 \$2215 \$1412 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$753 b2_r5_b_not \$2215 \$1195 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$754 \$2615 \$2217 b2_r5_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$755 \$1194 \$2070 \$2615 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$756 \$2616 \$2070 \$1195 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$757 b2_r5_b \$2217 \$2616 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$758 \$1194 \$2215 b2_r5_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$759 \$2095 a5|b0_p5|b1_p5|b3_p5|b4_p5|b5_p5|b6_p5|b7_p5 b2_c5_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$760 \$1420 \$2162 \$2095 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$761 \$2619 \$2163 \$1420 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$762 \$2096 \$2072 \$2619 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$763 \$2620 \$2072 \$2095 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$764 \$1421 \$2163 \$2620 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$765 \$2096 \$2162 \$1421 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$766 b3_r5_b_not \$2162 \$1202 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$767 \$2621 \$2163 b3_r5_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$768 \$1201 \$2072 \$2621 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$769 \$2622 \$2072 \$1202 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$770 b3_r5_b \$2163 \$2622 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$771 \$1201 \$2162 b3_r5_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$772 \$2100 b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b4|b4_q7 b2_c5_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$773 \$2623
+ b2_q0_not|b2_q1_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b4_not|b4_q7_not
+ \$2100 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$774 \$2102
+ a5_not|b0_p5_not|b1_p5_not|b2_p5_not|b3_p5_not|b5_p5_not|b6_p5_not|b7_p5_not
+ \$2623 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$775 \$2624
+ a5_not|b0_p5_not|b1_p5_not|b2_p5_not|b3_p5_not|b5_p5_not|b6_p5_not|b7_p5_not
+ b2_c5_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$776 \$2101
+ b2_q0_not|b2_q1_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b4_not|b4_q7_not
+ \$2624 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$777 \$2102 b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b4|b4_q7 \$2101 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$778 \$1429 \$2169 \$2100 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$779 \$2625 \$2224 \$1429 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$780 \$2101 \$2074 \$2625 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$781 \$2626 \$2074 \$2100 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$782 \$1430 \$2224 \$2626 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$783 \$2101 \$2169 \$1430 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$784 b4_r5_b_not \$2169 \$1206 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$785 \$2627 \$2224 b4_r5_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$786 \$1205 \$2074 \$2627 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$787 \$2628 \$2074 \$1206 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$788 b4_r5_b \$2224 \$2628 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$789 \$1205 \$2169 b4_r5_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$790 \$2106 b5|b5_q0|b5_q1|b5_q2|b5_q3|b5_q4|b5_q5|b5_q6|b5_q7 \$2105 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$791 \$2629
+ b5_not|b5_q0_not|b5_q1_not|b5_q2_not|b5_q3_not|b5_q4_not|b5_q5_not|b5_q6_not|b5_q7_not
+ \$2106 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$792 b5_c5
+ a5_not|b0_p5_not|b1_p5_not|b2_p5_not|b3_p5_not|b5_p5_not|b6_p5_not|b7_p5_not
+ \$2629 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$793 \$2630
+ a5_not|b0_p5_not|b1_p5_not|b2_p5_not|b3_p5_not|b5_p5_not|b6_p5_not|b7_p5_not
+ \$2105 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$794 \$2107
+ b5_not|b5_q0_not|b5_q1_not|b5_q2_not|b5_q3_not|b5_q4_not|b5_q5_not|b5_q6_not|b5_q7_not
+ \$2630 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$795 b5_c5 b5|b5_q0|b5_q1|b5_q2|b5_q3|b5_q4|b5_q5|b5_q6|b5_q7 \$2107 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$796 \$1438 \$2171 \$2106 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$797 \$2631 \$2229 \$1438 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$798 \$2107 \$2076 \$2631 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$799 \$2632 \$2076 \$2106 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$800 \$1439 \$2229 \$2632 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$801 \$2107 \$2171 \$1439 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$802 b5_r5_b_not \$2171 \$1210 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$803 \$2633 \$2229 b5_r5_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$804 \$1209 \$2076 \$2633 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$805 \$2634 \$2076 \$1210 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$806 b5_r5_b \$2229 \$2634 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$807 \$1209 \$2171 b5_r5_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$808 \$2111 b6|b6_q0|b6_q1|b6_q2|b6_q3|b6_q4|b6_q5|b6_q6|b6_q7 b6_c5_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$809 \$2111 a5|b0_p5|b1_p5|b3_p5|b4_p5|b5_p5|b6_p5|b7_p5 b6_c5_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$810 \$2635
+ b6_not|b6_q0_not|b6_q1_not|b6_q2_not|b6_q3_not|b6_q4_not|b6_q5_not|b6_q6_not|b6_q7_not
+ \$2111 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$811 b6_c5
+ a5_not|b0_p5_not|b1_p5_not|b2_p5_not|b3_p5_not|b5_p5_not|b6_p5_not|b7_p5_not
+ \$2635 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$812 \$2636
+ a5_not|b0_p5_not|b1_p5_not|b2_p5_not|b3_p5_not|b5_p5_not|b6_p5_not|b7_p5_not
+ b6_c5_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$813 \$2112
+ b6_not|b6_q0_not|b6_q1_not|b6_q2_not|b6_q3_not|b6_q4_not|b6_q5_not|b6_q6_not|b6_q7_not
+ \$2636 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$814 b6_c5 b6|b6_q0|b6_q1|b6_q2|b6_q3|b6_q4|b6_q5|b6_q6|b6_q7 \$2112 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$815 \$1447 \$2173 \$2111 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$816 \$2637 \$2236 \$1447 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$817 \$2112 \$2078 \$2637 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$818 \$2638 \$2078 \$2111 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$819 \$1448 \$2236 \$2638 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$820 \$2112 \$2173 \$1448 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$821 b6_r5_b_not \$2173 \$1214 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$822 \$2639 \$2236 b6_r5_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$823 \$1213 \$2078 \$2639 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$824 \$2640 \$2078 \$1214 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$825 b6_r5_b \$2236 \$2640 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$826 \$1213 \$2173 b6_r5_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$827 \$2116 b1_q3|b7|b7_q0|b7_q1|b7_q2|b7_q4|b7_q5|b7_q6|b7_q7 \$2115 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$828 \$2641
+ b7_not|b7_q0_not|b7_q1_not|b7_q2_not|b7_q3_not|b7_q4_not|b7_q5_not|b7_q6_not|b7_q7_not
+ \$2116 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$829 b6_c5
+ a5_not|b0_p5_not|b1_p5_not|b2_p5_not|b3_p5_not|b5_p5_not|b6_p5_not|b7_p5_not
+ \$2641 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$830 \$2642
+ a5_not|b0_p5_not|b1_p5_not|b2_p5_not|b3_p5_not|b5_p5_not|b6_p5_not|b7_p5_not
+ \$2115 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$831 \$2117
+ b7_not|b7_q0_not|b7_q1_not|b7_q2_not|b7_q3_not|b7_q4_not|b7_q5_not|b7_q6_not|b7_q7_not
+ \$2642 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$832 b6_c5 b1_q3|b7|b7_q0|b7_q1|b7_q2|b7_q4|b7_q5|b7_q6|b7_q7 \$2117 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$833 \$1456 \$2175 \$2116 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$834 \$2643 \$2241 \$1456 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$835 \$2117 \$2080 \$2643 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$836 \$2644 \$2080 \$2116 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$837 \$1457 \$2241 \$2644 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$838 \$2117 \$2175 \$1457 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$839 \$2118 \$2175 \$1218 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$840 \$2645 \$2241 \$2118 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$841 \$1217 \$2080 \$2645 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$842 \$2646 \$2080 \$1218 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$843 \$2119 \$2241 \$2646 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$844 \$1217 \$2175 \$2119 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$845 b1_c5 a5|b0_p5|b1_p5|b3_p5|b4_p5|b5_p5|b6_p5|b7_p5 \$2083 vdd pfet_03v3
+ L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$846 \$2090 a5|b0_p5|b1_p5|b3_p5|b4_p5|b5_p5|b6_p5|b7_p5 b2_c5_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$847 \$2100 a5|b0_p5|b1_p5|b3_p5|b4_p5|b5_p5|b6_p5|b7_p5 b2_c5_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$848 \$2106 a5|b0_p5|b1_p5|b3_p5|b4_p5|b5_p5|b6_p5|b7_p5 \$2105 vdd pfet_03v3
+ L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$849 \$2116 a5|b0_p5|b1_p5|b3_p5|b4_p5|b5_p5|b6_p5|b7_p5 \$2115 vdd pfet_03v3
+ L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$850 b0_c6 a6|b0_p6|b1_p6|b3_p6|b4_p6|b5_p6|b6_p6|b7_p6 \$2086 vdd pfet_03v3
+ L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$851 b3_c5 a5|b0_p5|b1_p5|b3_p5|b4_p5|b5_p5|b6_p5|b7_p5 \$2096 vdd pfet_03v3
+ L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$852 \$1420 \$2164 \$2095 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$853 b3_r5_b_not \$2164 \$1202 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$854 \$1429 \$2170 \$2100 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$855 \$1438 \$2172 \$2106 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$856 b6_c5 a5|b0_p5|b1_p5|b3_p5|b4_p5|b5_p5|b6_p5|b7_p5 \$2112 vdd pfet_03v3
+ L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$857 \$1447 \$2174 \$2111 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$858 \$1456 \$2176 \$2116 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$859 \$1402 \$2209 \$2085 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$860 b0_r6_b_not \$2209 \$1191 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$861 b2_c5 a5|b0_p5|b1_p5|b3_p5|b4_p5|b5_p5|b6_p5|b7_p5 \$2091 vdd pfet_03v3
+ L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$862 \$1411 \$2216 \$2090 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$863 b2_r5_b_not \$2216 \$1195 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$864 \$2096 \$2164 \$1421 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$865 \$1201 \$2164 b3_r5_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$866 \$2102 a5|b0_p5|b1_p5|b3_p5|b4_p5|b5_p5|b6_p5|b7_p5 \$2101 vdd pfet_03v3
+ L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$867 \$2101 \$2170 \$1430 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$868 b4_r5_b_not \$2170 \$1206 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$869 b5_c5 a5|b0_p5|b1_p5|b3_p5|b4_p5|b5_p5|b6_p5|b7_p5 \$2107 vdd pfet_03v3
+ L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$870 \$2107 \$2172 \$1439 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$871 b5_r5_b_not \$2172 \$1210 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$872 \$2112 \$2174 \$1448 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$873 b6_r5_b_not \$2174 \$1214 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$874 b6_c5 a5|b0_p5|b1_p5|b3_p5|b4_p5|b5_p5|b6_p5|b7_p5 \$2117 vdd pfet_03v3
+ L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$875 \$2117 \$2176 \$1457 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$876 \$2118 \$2176 \$1218 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$877 \$2086 \$2209 \$1403 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$878 \$1190 \$2209 b0_r6_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$879 \$2091 \$2216 \$1412 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$880 \$1194 \$2216 b2_r5_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$881 \$3189 \$3057 \$2221 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$882 \$2220 \$3058 \$3189 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$883 \$2221 \$3058 \$3191 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$884 \$3190 \$3057 \$3118 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$885 \$3342 \$3058 \$3190 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$886 \$3118 \$3058 \$3036 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$887 \$3119 b3_r4_b_not \$3036 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$888 \$3190 b3_r4_b \$3119 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$889 \$3036 b3_r4_b \$3120 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$890 \$3121 \$3120 \$3191 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$891 \$3189 \$3119 \$3121 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$892 \$3191 \$3119 \$3122 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$893 \$1205 \$2170 b4_r5_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$894 \$3195 b4_r4_b_not \$3037 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$895 \$3037 b4_r4_b \$3124 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$896 \$3196 \$3124 \$3194 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$897 \$3194 \$3195 \$3125 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$898 \$1209 \$2172 b5_r5_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$899 \$3200 b5_r4_b_not \$3038 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$900 \$3038 b5_r4_b \$3127 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$901 \$3201 \$3127 \$3199 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$902 \$3199 \$3200 \$3128 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$903 \$1213 \$2174 b6_r5_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$904 \$3205 b6_r4_b_not \$3039 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$905 \$3039 b6_r4_b \$3130 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$906 \$3206 \$3130 \$3204 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$907 \$3204 \$3205 \$3131 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$908 \$1217 \$2176 \$2119 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$909 \$3210 \$3085 \$3040 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$910 \$3040 \$3086 \$3133 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$911 p11 \$3133 \$3209 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$912 \$3209 \$3210 p11_not vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$913 \$3178 b0_r5_b_not \$3034 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$914 \$3176 b0_r5_b \$3178 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$915 \$3034 b0_r5_b \$3179 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$916 \$3180 \$3179 \$3177 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$917 \$3175 \$3178 \$3180 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$918 \$3177 \$3178 \$3181 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$919 \$3185 b2_r4_b_not \$3035 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$920 \$3183 b2_r4_b \$3185 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$921 \$3035 b2_r4_b \$3186 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$922 \$3187 \$3186 \$3184 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$923 \$3182 \$3185 \$3187 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$924 \$3184 \$3185 \$3188 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$925 \$3120 b3_r4_b_not \$3190 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$926 \$3122 \$3120 \$3189 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$927 \$3192 \$3062 \$2168 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$928 \$2168 \$3064 \$3194 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$929 \$3193 \$3062 \$3123 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$930 \$3123 \$3064 \$3037 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$931 \$3193 b4_r4_b \$3195 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$932 \$3192 \$3195 \$3196 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$933 \$3197 \$3068 \$2228 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$934 \$2228 \$3070 \$3199 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$935 \$3198 \$3068 \$3126 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$936 \$3126 \$3070 \$3038 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$937 \$3198 b5_r4_b \$3200 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$938 \$3197 \$3200 \$3201 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$939 \$3202 \$3075 \$2233 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$940 \$2233 \$3077 \$3204 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$941 \$3203 \$3075 \$3129 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$942 \$3129 \$3077 \$3039 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$943 \$3203 b6_r4_b \$3205 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$944 \$3202 \$3205 \$3206 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$945 \$3207 \$3081 \$2240 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$946 \$2240 \$3083 \$3209 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$947 \$3208 \$3081 \$3132 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$948 \$3132 \$3083 \$3040 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$949 \$3208 \$3086 \$3210 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$950 \$3207 \$3210 p11 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$951 \$3115 b1|b1_q0|b1_q1|b1_q2|b1_q3|b1_q4|b1_q5|b1_q6|b1_q7 b1_c4_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$952 \$3570
+ b1_not|b1_q0_not|b1_q1_not|b1_q2_not|b1_q3_not|b1_q4_not|b1_q5_not|b1_q6_not|b1_q7_not
+ \$3115 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$953 b1_c4
+ a4_not|b0_p4_not|b1_p4_not|b2_p4_not|b3_p4_not|b5_p4_not|b6_p4_not|b7_p4_not
+ \$3570 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$954 \$3571
+ a4_not|b0_p4_not|b1_p4_not|b2_p4_not|b3_p4_not|b5_p4_not|b6_p4_not|b7_p4_not
+ b1_c4_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$955 \$3043
+ b1_not|b1_q0_not|b1_q1_not|b1_q2_not|b1_q3_not|b1_q4_not|b1_q5_not|b1_q6_not|b1_q7_not
+ \$3571 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$956 b1_c4 b1|b1_q0|b1_q1|b1_q2|b1_q3|b1_q4|b1_q5|b1_q6|b1_q7 \$3043 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$957 \$3175 \$3045 \$3115 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$958 \$3043 \$3047 \$3175 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$959 \$3177 \$3045 \$3043 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$960 \$3115 \$3047 \$3177 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$961 \$3176 \$3045 \$3116 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$962 \$3328 \$3047 \$3176 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$963 \$3034 \$3045 \$3328 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$964 \$3116 \$3047 \$3034 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$965 \$3179 b0_r5_b_not \$3176 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$966 \$3181 \$3179 \$3175 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$967 \$3182 \$3051 \$2214 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$968 \$2213 \$3053 \$3182 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$969 \$3184 \$3051 \$2213 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$970 \$2214 \$3053 \$3184 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$971 \$3183 \$3051 \$3117 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$972 \$3335 \$3053 \$3183 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$973 \$3035 \$3051 \$3335 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$974 \$3117 \$3053 \$3035 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P AD=0.70395P
+ PS=3.51U PD=3.61U
M$975 \$3186 b2_r4_b_not \$3183 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$976 \$3188 \$3186 \$3182 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$977 \$3057
+ b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b3|b3_q0|b3_q1|b3_q2|b3_q3|b3_q4|b3_q5|b3_q6|b3_q7
+ b2_c4_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$978 \$3580
+ b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b3_not|b3_q0_not|b3_q1_not|b3_q2_not|b3_q3_not|b3_q4_not|b3_q5_not|b3_q6_not|b3_q7_not
+ \$3057 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$979 b2_c4
+ a4_not|b0_p4_not|b1_p4_not|b2_p4_not|b3_p4_not|b5_p4_not|b6_p4_not|b7_p4_not
+ \$3580 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$980 \$3581
+ a4_not|b0_p4_not|b1_p4_not|b2_p4_not|b3_p4_not|b5_p4_not|b6_p4_not|b7_p4_not
+ b2_c4_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$981 \$3058
+ b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b3_not|b3_q0_not|b3_q1_not|b3_q2_not|b3_q3_not|b3_q4_not|b3_q5_not|b3_q6_not|b3_q7_not
+ \$3581 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$982 b2_c4
+ b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b3|b3_q0|b3_q1|b3_q2|b3_q3|b3_q4|b3_q5|b3_q6|b3_q7
+ \$3058 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$983 \$3191 \$3057 \$2220 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$984 \$3036 \$3057 \$3342 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$985 \$2375 \$3189 \$3057 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$986 \$3582 \$3191 \$2375 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$987 \$3058 \$3036 \$3582 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$988 \$3583 \$3036 \$3057 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$989 \$2376 \$3191 \$3583 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$990 \$3058 \$3189 \$2376 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$991 b3_r4_b_not \$3189 \$2166 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$992 \$3584 \$3191 b3_r4_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$993 \$2165 \$3036 \$3584 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$994 \$3585 \$3036 \$2166 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$995 b3_r4_b \$3191 \$3585 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$996 \$2165 \$3189 b3_r4_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$997 \$2167 \$3064 \$3192 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$998 \$3194 \$3062 \$2167 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$999 \$3349 \$3064 \$3193 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$1000 \$3037 \$3062 \$3349 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1001 \$3124 b4_r4_b_not \$3193 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1002 \$3125 \$3124 \$3192 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1003 \$2227 \$3070 \$3197 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1004 \$3199 \$3068 \$2227 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1005 \$3356 \$3070 \$3198 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1006 \$3038 \$3068 \$3356 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1007 \$3127 b5_r4_b_not \$3198 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1008 \$3128 \$3127 \$3197 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1009 \$2232 \$3077 \$3202 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1010 \$3204 \$3075 \$2232 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1011 \$3364 \$3077 \$3203 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1012 \$3039 \$3075 \$3364 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1013 \$3130 b6_r4_b_not \$3203 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1014 \$3131 \$3130 \$3202 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1015 \$2239 \$3083 \$3207 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1016 \$3209 \$3081 \$2239 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1017 \$3371 \$3083 \$3208 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1018 \$3040 \$3081 \$3371 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1019 \$3133 \$3085 \$3208 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1020 p11_not \$3133 \$3207 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1021 \$3115 a4|b0_p4|b1_p4|b2_p4|b3_p4|b4_p4|b5_p4|b6_p4|b7_p4 b1_c4_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1022 b1_c4 a4|b0_p4|b1_p4|b2_p4|b3_p4|b4_p4|b5_p4|b6_p4|b7_p4 \$3043 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1023 \$3045 b0|b0_q0|b0_q1|b0_q2|b0_q3|b0_q4|b0_q5|b0_q6|b0_q7 b0_c5_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1024 \$3045 a5|b0_p5|b1_p5|b3_p5|b4_p5|b5_p5|b6_p5|b7_p5 b0_c5_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1025 \$3572
+ b0_not|b0_q0_not|b0_q1_not|b0_q3_not|b0_q4_not|b0_q5_not|b0_q6_not|b0_q7_not|b1_q2_not
+ \$3045 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1026 b0_c5
+ a5_not|b0_p5_not|b1_p5_not|b2_p5_not|b3_p5_not|b5_p5_not|b6_p5_not|b7_p5_not
+ \$3572 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1027 \$3573
+ a5_not|b0_p5_not|b1_p5_not|b2_p5_not|b3_p5_not|b5_p5_not|b6_p5_not|b7_p5_not
+ b0_c5_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1028 \$3047
+ b0_not|b0_q0_not|b0_q1_not|b0_q3_not|b0_q4_not|b0_q5_not|b0_q6_not|b0_q7_not|b1_q2_not
+ \$3573 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1029 b0_c5 b0|b0_q0|b0_q1|b0_q2|b0_q3|b0_q4|b0_q5|b0_q6|b0_q7 \$3047 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1030 b0_c5 a5|b0_p5|b1_p5|b3_p5|b4_p5|b5_p5|b6_p5|b7_p5 \$3047 vdd pfet_03v3
+ L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1031 \$2360 \$3176 \$3045 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1032 \$2360 \$3175 \$3045 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1033 \$3613 \$3177 \$2360 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1034 \$3047 \$3034 \$3613 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1035 \$3614 \$3034 \$3045 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1036 \$2361 \$3177 \$3614 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1037 \$3047 \$3175 \$2361 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1038 b0_r5_b_not \$3175 \$2212 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1039 b0_r5_b_not \$3176 \$2212 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1040 \$3574 \$3177 b0_r5_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1041 \$2211 \$3034 \$3574 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1042 \$3575 \$3034 \$2212 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1043 b0_r5_b \$3177 \$3575 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1044 \$2211 \$3175 b0_r5_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1045 \$3051 b2|b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7 b2_c4_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1046 \$3051 a4|b0_p4|b1_p4|b2_p4|b3_p4|b4_p4|b5_p4|b6_p4|b7_p4 b2_c4_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1047 \$3576
+ b2_not|b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not
+ \$3051 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1048 b2_c4
+ a4_not|b0_p4_not|b1_p4_not|b2_p4_not|b3_p4_not|b5_p4_not|b6_p4_not|b7_p4_not
+ \$3576 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1049 \$3577
+ a4_not|b0_p4_not|b1_p4_not|b2_p4_not|b3_p4_not|b5_p4_not|b6_p4_not|b7_p4_not
+ b2_c4_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1050 \$3053
+ b2_not|b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not
+ \$3577 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1051 b2_c4 b2|b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7 \$3053 vdd pfet_03v3
+ L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1052 \$2368 \$3182 \$3051 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1053 \$2368 \$3183 \$3051 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1054 \$3617 \$3184 \$2368 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1055 \$3053 \$3035 \$3617 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1056 \$3618 \$3035 \$3051 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1057 \$2369 \$3184 \$3618 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1058 \$3053 \$3182 \$2369 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1059 b2_r4_b_not \$3183 \$2219 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1060 b2_r4_b_not \$3182 \$2219 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1061 \$3578 \$3184 b2_r4_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1062 \$2218 \$3035 \$3578 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1063 \$3579 \$3035 \$2219 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1064 b2_r4_b \$3184 \$3579 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1065 \$2218 \$3182 b2_r4_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1066 \$3057 a4|b0_p4|b1_p4|b2_p4|b3_p4|b4_p4|b5_p4|b6_p4|b7_p4 b2_c4_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1067 b2_c4 a4|b0_p4|b1_p4|b2_p4|b3_p4|b4_p4|b5_p4|b6_p4|b7_p4 \$3058 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1068 \$2375 \$3190 \$3057 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1069 \$3058 \$3190 \$2376 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1070 b3_r4_b_not \$3190 \$2166 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1071 \$2165 \$3190 b3_r4_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1072 \$3062 b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b4|b4_q7 b2_c4_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1073 \$3062 a4|b0_p4|b1_p4|b2_p4|b3_p4|b4_p4|b5_p4|b6_p4|b7_p4 b2_c4_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1074 \$3586
+ b2_q0_not|b2_q1_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b4_not|b4_q7_not
+ \$3062 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1075 b2_c4
+ a4_not|b0_p4_not|b1_p4_not|b2_p4_not|b3_p4_not|b5_p4_not|b6_p4_not|b7_p4_not
+ \$3586 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1076 \$3587
+ a4_not|b0_p4_not|b1_p4_not|b2_p4_not|b3_p4_not|b5_p4_not|b6_p4_not|b7_p4_not
+ b2_c4_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1077 \$3064
+ b2_q0_not|b2_q1_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b4_not|b4_q7_not
+ \$3587 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1078 b2_c4 b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b4|b4_q7 \$3064 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1079 \$2383 \$3192 \$3062 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1080 \$2383 \$3193 \$3062 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1081 \$3588 \$3194 \$2383 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1082 \$3064 \$3037 \$3588 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1083 \$3589 \$3037 \$3062 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1084 \$2384 \$3194 \$3589 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1085 \$3064 \$3192 \$2384 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1086 b4_r4_b_not \$3193 \$2226 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1087 b4_r4_b_not \$3192 \$2226 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1088 \$3590 \$3194 b4_r4_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1089 \$2225 \$3037 \$3590 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1090 \$3591 \$3037 \$2226 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1091 b4_r4_b \$3194 \$3591 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1092 \$2225 \$3193 b4_r4_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1093 \$2225 \$3192 b4_r4_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1094 \$3068 b5|b5_q0|b5_q1|b5_q2|b5_q3|b5_q4|b5_q5|b5_q6|b5_q7 \$3067 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1095 \$3068 a4|b0_p4|b1_p4|b2_p4|b3_p4|b4_p4|b5_p4|b6_p4|b7_p4 \$3067 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1096 \$3592
+ b5_not|b5_q0_not|b5_q1_not|b5_q2_not|b5_q3_not|b5_q4_not|b5_q5_not|b5_q6_not|b5_q7_not
+ \$3068 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1097 \$3071
+ a4_not|b0_p4_not|b1_p4_not|b2_p4_not|b3_p4_not|b5_p4_not|b6_p4_not|b7_p4_not
+ \$3592 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1098 \$3593
+ a4_not|b0_p4_not|b1_p4_not|b2_p4_not|b3_p4_not|b5_p4_not|b6_p4_not|b7_p4_not
+ \$3067 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1099 \$3070
+ b5_not|b5_q0_not|b5_q1_not|b5_q2_not|b5_q3_not|b5_q4_not|b5_q5_not|b5_q6_not|b5_q7_not
+ \$3593 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1100 \$3071 b5|b5_q0|b5_q1|b5_q2|b5_q3|b5_q4|b5_q5|b5_q6|b5_q7 \$3070 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1101 \$2391 \$3198 \$3068 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1102 \$2391 \$3197 \$3068 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1103 \$3594 \$3199 \$2391 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1104 \$3070 \$3038 \$3594 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1105 \$3595 \$3038 \$3068 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1106 \$2392 \$3199 \$3595 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1107 \$3070 \$3197 \$2392 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1108 b5_r4_b_not \$3198 \$2231 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1109 b5_r4_b_not \$3197 \$2231 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1110 \$3596 \$3199 b5_r4_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1111 \$2230 \$3038 \$3596 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1112 \$3597 \$3038 \$2231 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1113 b5_r4_b \$3199 \$3597 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1114 \$2230 \$3197 b5_r4_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1115 \$2230 \$3198 b5_r4_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1116 \$3075 b6|b6_q0|b6_q1|b6_q2|b6_q3|b6_q4|b6_q5|b6_q6|b6_q7 b6_c4_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1117 \$3075 a4|b0_p4|b1_p4|b2_p4|b3_p4|b4_p4|b5_p4|b6_p4|b7_p4 b6_c4_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1118 \$3598
+ b6_not|b6_q0_not|b6_q1_not|b6_q2_not|b6_q3_not|b6_q4_not|b6_q5_not|b6_q6_not|b6_q7_not
+ \$3075 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1119 b6_c4
+ a4_not|b0_p4_not|b1_p4_not|b2_p4_not|b3_p4_not|b5_p4_not|b6_p4_not|b7_p4_not
+ \$3598 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1120 \$3599
+ a4_not|b0_p4_not|b1_p4_not|b2_p4_not|b3_p4_not|b5_p4_not|b6_p4_not|b7_p4_not
+ b6_c4_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1121 \$3077
+ b6_not|b6_q0_not|b6_q1_not|b6_q2_not|b6_q3_not|b6_q4_not|b6_q5_not|b6_q6_not|b6_q7_not
+ \$3599 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1122 b6_c4 b6|b6_q0|b6_q1|b6_q2|b6_q3|b6_q4|b6_q5|b6_q6|b6_q7 \$3077 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1123 \$2398 \$3202 \$3075 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1124 \$2398 \$3203 \$3075 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1125 \$3600 \$3204 \$2398 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1126 \$3077 \$3039 \$3600 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1127 \$3601 \$3039 \$3075 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1128 \$2399 \$3204 \$3601 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1129 \$3077 \$3202 \$2399 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1130 b6_r4_b_not \$3203 \$2238 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1131 b6_r4_b_not \$3202 \$2238 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1132 \$3602 \$3204 b6_r4_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1133 \$2237 \$3039 \$3602 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1134 \$3603 \$3039 \$2238 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1135 b6_r4_b \$3204 \$3603 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1136 \$2237 \$3203 b6_r4_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1137 \$2237 \$3202 b6_r4_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1138 \$3081 b1_q3|b7|b7_q0|b7_q1|b7_q2|b7_q4|b7_q5|b7_q6|b7_q7 \$3080 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1139 \$3081 a4|b0_p4|b1_p4|b2_p4|b3_p4|b4_p4|b5_p4|b6_p4|b7_p4 \$3080 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1140 \$3604
+ b7_not|b7_q0_not|b7_q1_not|b7_q2_not|b7_q3_not|b7_q4_not|b7_q5_not|b7_q6_not|b7_q7_not
+ \$3081 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1141 \$3084
+ a4_not|b0_p4_not|b1_p4_not|b2_p4_not|b3_p4_not|b5_p4_not|b6_p4_not|b7_p4_not
+ \$3604 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1142 \$3605
+ a4_not|b0_p4_not|b1_p4_not|b2_p4_not|b3_p4_not|b5_p4_not|b6_p4_not|b7_p4_not
+ \$3080 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1143 \$3083
+ b7_not|b7_q0_not|b7_q1_not|b7_q2_not|b7_q3_not|b7_q4_not|b7_q5_not|b7_q6_not|b7_q7_not
+ \$3605 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1144 \$3084 b1_q3|b7|b7_q0|b7_q1|b7_q2|b7_q4|b7_q5|b7_q6|b7_q7 \$3083 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1145 \$2406 \$3208 \$3081 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1146 \$2406 \$3207 \$3081 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1147 \$3606 \$3209 \$2406 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1148 \$3083 \$3040 \$3606 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1149 \$3607 \$3040 \$3081 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1150 \$2407 \$3209 \$3607 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1151 \$3083 \$3207 \$2407 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1152 \$3085 \$3207 \$2243 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1153 \$3085 \$3208 \$2243 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1154 \$3608 \$3209 \$3085 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1155 \$2242 \$3040 \$3608 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1156 \$3609 \$3040 \$2243 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1157 \$3086 \$3209 \$3609 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1158 \$2242 \$3208 \$3086 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1159 \$2242 \$3207 \$3086 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1160 \$3047 \$3176 \$2361 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1161 \$2211 \$3176 b0_r5_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1162 b2_c4 a4|b0_p4|b1_p4|b2_p4|b3_p4|b4_p4|b5_p4|b6_p4|b7_p4 \$3053 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1163 \$3053 \$3183 \$2369 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1164 \$2218 \$3183 b2_r4_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1165 \$4087 \$4051 \$3188 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1166 \$3187 \$4052 \$4087 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1167 \$3188 \$4052 \$4159 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1168 \$4088 \$4051 \$4089 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1169 \$4309 \$4052 \$4088 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1170 \$4089 \$4052 \$3620 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1171 \$4090 b3_r3_b_not \$3620 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1172 \$4088 b3_r3_b \$4090 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1173 \$3620 b3_r3_b \$4091 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1174 \$4092 \$4091 \$4159 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1175 \$4087 \$4090 \$4092 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1176 \$4159 \$4090 \$4093 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1177 b2_c4 a4|b0_p4|b1_p4|b2_p4|b3_p4|b4_p4|b5_p4|b6_p4|b7_p4 \$3064 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1178 \$3122 \$4057 \$4160 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1179 \$4096 \$4057 \$3622 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1180 \$3064 \$3193 \$2384 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1181 \$3071 a4|b0_p4|b1_p4|b2_p4|b3_p4|b4_p4|b5_p4|b6_p4|b7_p4 \$3070 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1182 \$3125 \$4062 \$4165 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1183 \$4099 \$4062 \$3624 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1184 \$3070 \$3198 \$2392 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1185 b6_c4 a4|b0_p4|b1_p4|b2_p4|b3_p4|b4_p4|b5_p4|b6_p4|b7_p4 \$3077 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1186 \$3128 \$4067 \$4170 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1187 \$4102 \$4067 \$3626 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1188 \$3077 \$3203 \$2399 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1189 \$3084 a4|b0_p4|b1_p4|b2_p4|b3_p4|b4_p4|b5_p4|b6_p4|b7_p4 \$3083 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1190 \$3131 \$4072 \$4175 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1191 \$4105 \$4072 \$3628 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1192 \$3083 \$3208 \$2407 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1193 \$4038 \$4042 \$4147 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1194 \$4085 \$4042 \$3612 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1195 \$3181 \$4047 \$4154 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1196 \$4086 \$4047 \$3616 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1197 \$4094 \$4056 \$3122 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1198 \$3121 \$4057 \$4094 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1199 \$4095 \$4056 \$4096 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1200 \$4317 \$4057 \$4095 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1201 \$4097 \$4061 \$3125 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1202 \$3196 \$4062 \$4097 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1203 \$4098 \$4061 \$4099 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1204 \$4325 \$4062 \$4098 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1205 \$4100 \$4066 \$3128 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1206 \$3201 \$4067 \$4100 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1207 \$4101 \$4066 \$4102 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1208 \$4332 \$4067 \$4101 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1209 \$4103 \$4071 \$3131 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1210 \$3206 \$4072 \$4103 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1211 \$4104 \$4071 \$4105 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1212 \$4340 \$4072 \$4104 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1213 \$4145 \$4041 \$4038 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1214 \$4039 \$4042 \$4145 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1215 \$4146 \$4041 \$4085 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1216 \$4293 \$4042 \$4146 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1217 \$4148 b0_r4_b_not \$3612 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1218 \$3612 b0_r4_b \$4149 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1219 \$4150 \$4149 \$4147 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1220 \$4147 \$4148 \$4151 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1221 \$4152 \$4046 \$3181 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1222 \$3180 \$4047 \$4152 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1223 \$4153 \$4046 \$4086 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1224 \$4301 \$4047 \$4153 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1225 \$4155 b2_r3_b_not \$3616 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1226 \$3616 b2_r3_b \$4156 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1227 \$4157 \$4156 \$4154 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1228 \$4154 \$4155 \$4158 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1229 \$4159 \$4051 \$3187 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1230 \$3620 \$4051 \$4309 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1231 \$4091 b3_r3_b_not \$4088 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1232 \$4093 \$4091 \$4087 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1233 \$4161 b4_r3_b_not \$3622 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1234 \$4095 b4_r3_b \$4161 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1235 \$3622 b4_r3_b \$4162 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1236 \$4163 \$4162 \$4160 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1237 \$4094 \$4161 \$4163 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1238 \$4160 \$4161 \$4164 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1239 \$4166 b5_r3_b_not \$3624 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1240 \$4098 b5_r3_b \$4166 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1241 \$3624 b5_r3_b \$4167 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1242 \$4168 \$4167 \$4165 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1243 \$4097 \$4166 \$4168 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1244 \$4165 \$4166 \$4169 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1245 \$4171 b6_r3_b_not \$3626 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1246 \$4101 b6_r3_b \$4171 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1247 \$3626 b6_r3_b \$4172 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1248 \$4173 \$4172 \$4170 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1249 \$4100 \$4171 \$4173 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1250 \$4170 \$4171 \$4174 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1251 \$4176 \$4073 \$3628 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1252 \$4104 \$4074 \$4176 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1253 \$3628 \$4074 \$4177 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1254 p10 \$4177 \$4175 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$1255 \$4103 \$4176 p10 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$1256 \$4175 \$4176 p10_not vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1257 \$4038 b1|b1_q0|b1_q1|b1_q2|b1_q3|b1_q4|b1_q5|b1_q6|b1_q7 b1_c3_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1258 \$4537
+ b1_not|b1_q0_not|b1_q1_not|b1_q2_not|b1_q3_not|b1_q4_not|b1_q5_not|b1_q6_not|b1_q7_not
+ \$4038 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1259 b1_c3
+ a3_not|b0_p3_not|b1_p3_not|b2_p3_not|b3_p3_not|b5_p3_not|b6_p3_not|b7_p3_not
+ \$4537 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1260 \$4538
+ a3_not|b0_p3_not|b1_p3_not|b2_p3_not|b3_p3_not|b5_p3_not|b6_p3_not|b7_p3_not
+ b1_c3_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1261 \$4039
+ b1_not|b1_q0_not|b1_q1_not|b1_q2_not|b1_q3_not|b1_q4_not|b1_q5_not|b1_q6_not|b1_q7_not
+ \$4538 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1262 b1_c3 b1|b1_q0|b1_q1|b1_q2|b1_q3|b1_q4|b1_q5|b1_q6|b1_q7 \$4039 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1263 \$4041 b0|b0_q0|b0_q1|b0_q2|b0_q3|b0_q4|b0_q5|b0_q6|b0_q7 b0_c4_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1264 \$4539
+ b0_not|b0_q0_not|b0_q1_not|b0_q3_not|b0_q4_not|b0_q5_not|b0_q6_not|b0_q7_not|b1_q2_not
+ \$4041 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1265 b0_c4
+ a4_not|b0_p4_not|b1_p4_not|b2_p4_not|b3_p4_not|b5_p4_not|b6_p4_not|b7_p4_not
+ \$4539 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1266 \$4540
+ a4_not|b0_p4_not|b1_p4_not|b2_p4_not|b3_p4_not|b5_p4_not|b6_p4_not|b7_p4_not
+ b0_c4_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1267 \$4042
+ b0_not|b0_q0_not|b0_q1_not|b0_q3_not|b0_q4_not|b0_q5_not|b0_q6_not|b0_q7_not|b1_q2_not
+ \$4540 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1268 b0_c4 b0|b0_q0|b0_q1|b0_q2|b0_q3|b0_q4|b0_q5|b0_q6|b0_q7 \$4042 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1269 \$4147 \$4041 \$4039 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1270 \$3612 \$4041 \$4293 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1271 \$4146 b0_r4_b \$4148 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1272 \$4149 b0_r4_b_not \$4146 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1273 \$4145 \$4148 \$4150 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1274 \$4151 \$4149 \$4145 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1275 \$4046 b2|b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7 b2_c2_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1276 \$4545
+ b2_not|b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not
+ \$4046 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1277 b2_c2
+ a3_not|b0_p3_not|b1_p3_not|b2_p3_not|b3_p3_not|b5_p3_not|b6_p3_not|b7_p3_not
+ \$4545 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1278 \$4546
+ a3_not|b0_p3_not|b1_p3_not|b2_p3_not|b3_p3_not|b5_p3_not|b6_p3_not|b7_p3_not
+ b2_c2_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1279 \$4047
+ b2_not|b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not
+ \$4546 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1280 b2_c2 b2|b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7 \$4047 vdd pfet_03v3
+ L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1281 \$4154 \$4046 \$3180 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1282 \$3616 \$4046 \$4301 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1283 \$4153 b2_r3_b \$4155 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1284 \$4156 b2_r3_b_not \$4153 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1285 \$4152 \$4155 \$4157 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1286 \$4158 \$4156 \$4152 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1287 \$4051
+ b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b3|b3_q0|b3_q1|b3_q2|b3_q3|b3_q4|b3_q5|b3_q6|b3_q7
+ b3_c2_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1288 \$4551
+ b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b3_not|b3_q0_not|b3_q1_not|b3_q2_not|b3_q3_not|b3_q4_not|b3_q5_not|b3_q6_not|b3_q7_not
+ \$4051 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1289 b3_c2
+ a3_not|b0_p3_not|b1_p3_not|b2_p3_not|b3_p3_not|b5_p3_not|b6_p3_not|b7_p3_not
+ \$4551 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1290 \$4552
+ a3_not|b0_p3_not|b1_p3_not|b2_p3_not|b3_p3_not|b5_p3_not|b6_p3_not|b7_p3_not
+ b3_c2_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1291 \$4052
+ b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b3_not|b3_q0_not|b3_q1_not|b3_q2_not|b3_q3_not|b3_q4_not|b3_q5_not|b3_q6_not|b3_q7_not
+ \$4552 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1292 b3_c2
+ b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b3|b3_q0|b3_q1|b3_q2|b3_q3|b3_q4|b3_q5|b3_q6|b3_q7
+ \$4052 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1293 \$3118 \$4087 \$4051 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1294 \$4553 \$4159 \$3118 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1295 \$4052 \$3620 \$4553 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1296 \$4554 \$3620 \$4051 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1297 \$3342 \$4159 \$4554 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1298 \$4052 \$4087 \$3342 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1299 b3_r3_b_not \$4087 \$3120 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1300 \$4555 \$4159 b3_r3_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1301 \$3119 \$3620 \$4555 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1302 \$4556 \$3620 \$3120 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1303 b3_r3_b \$4159 \$4556 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1304 \$3119 \$4087 b3_r3_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1305 \$4160 \$4056 \$3121 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1306 \$3622 \$4056 \$4317 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1307 \$3123 \$4094 \$4056 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1308 \$4559 \$4160 \$3123 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1309 \$4057 \$3622 \$4559 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1310 \$4560 \$3622 \$4056 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1311 \$3349 \$4160 \$4560 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1312 \$4057 \$4094 \$3349 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1313 \$4162 b4_r3_b_not \$4095 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1314 \$4164 \$4162 \$4094 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1315 \$4165 \$4061 \$3196 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1316 \$3624 \$4061 \$4325 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1317 \$3126 \$4097 \$4061 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1318 \$4565 \$4165 \$3126 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1319 \$4062 \$3624 \$4565 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1320 \$4566 \$3624 \$4061 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1321 \$3356 \$4165 \$4566 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1322 \$4062 \$4097 \$3356 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1323 \$4167 b5_r3_b_not \$4098 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1324 \$4169 \$4167 \$4097 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1325 \$4066 b6|b6_q0|b6_q1|b6_q2|b6_q3|b6_q4|b6_q5|b6_q6|b6_q7
+ b6_c2_not|b6_c3_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1326 \$4569
+ b6_not|b6_q0_not|b6_q1_not|b6_q2_not|b6_q3_not|b6_q4_not|b6_q5_not|b6_q6_not|b6_q7_not
+ \$4066 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1327 b6_c2|b6_c3
+ a3_not|b0_p3_not|b1_p3_not|b2_p3_not|b3_p3_not|b5_p3_not|b6_p3_not|b7_p3_not
+ \$4569 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1328 \$4570
+ a3_not|b0_p3_not|b1_p3_not|b2_p3_not|b3_p3_not|b5_p3_not|b6_p3_not|b7_p3_not
+ b6_c2_not|b6_c3_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1329 \$4067
+ b6_not|b6_q0_not|b6_q1_not|b6_q2_not|b6_q3_not|b6_q4_not|b6_q5_not|b6_q6_not|b6_q7_not
+ \$4570 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1330 b6_c2|b6_c3 b6|b6_q0|b6_q1|b6_q2|b6_q3|b6_q4|b6_q5|b6_q6|b6_q7 \$4067
+ vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1331 \$4170 \$4066 \$3201 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1332 \$3626 \$4066 \$4332 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1333 \$3129 \$4100 \$4066 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1334 \$4571 \$4170 \$3129 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1335 \$4067 \$3626 \$4571 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1336 \$4572 \$3626 \$4066 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1337 \$3364 \$4170 \$4572 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1338 \$4067 \$4100 \$3364 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1339 \$4172 b6_r3_b_not \$4101 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1340 \$4174 \$4172 \$4100 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1341 \$4071 b1_q3|b7|b7_q0|b7_q1|b7_q2|b7_q4|b7_q5|b7_q6|b7_q7 b6_c2_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1342 \$4575
+ b7_not|b7_q0_not|b7_q1_not|b7_q2_not|b7_q3_not|b7_q4_not|b7_q5_not|b7_q6_not|b7_q7_not
+ \$4071 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1343 b6_c2
+ a3_not|b0_p3_not|b1_p3_not|b2_p3_not|b3_p3_not|b5_p3_not|b6_p3_not|b7_p3_not
+ \$4575 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1344 \$4576
+ a3_not|b0_p3_not|b1_p3_not|b2_p3_not|b3_p3_not|b5_p3_not|b6_p3_not|b7_p3_not
+ b6_c2_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1345 \$4072
+ b7_not|b7_q0_not|b7_q1_not|b7_q2_not|b7_q3_not|b7_q4_not|b7_q5_not|b7_q6_not|b7_q7_not
+ \$4576 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1346 b6_c2 b1_q3|b7|b7_q0|b7_q1|b7_q2|b7_q4|b7_q5|b7_q6|b7_q7 \$4072 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1347 \$4175 \$4071 \$3206 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1348 \$3628 \$4071 \$4340 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1349 \$3132 \$4103 \$4071 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1350 \$4577 \$4175 \$3132 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1351 \$4072 \$3628 \$4577 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1352 \$4578 \$3628 \$4071 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1353 \$3371 \$4175 \$4578 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1354 \$4072 \$4103 \$3371 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1355 \$4177 \$4073 \$4104 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1356 p10_not \$4177 \$4103 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1357 \$4038 a3|b0_p3|b1_p3|b2_p3|b3_p3|b5_p3|b6_p3|b7_p3 b1_c3_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1358 b1_c3 a3|b0_p3|b1_p3|b2_p3|b3_p3|b5_p3|b6_p3|b7_p3 \$4039 vdd pfet_03v3
+ L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1359 \$4041 a4|b0_p4|b1_p4|b2_p4|b3_p4|b4_p4|b5_p4|b6_p4|b7_p4 b0_c4_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1360 b0_c4 a4|b0_p4|b1_p4|b2_p4|b3_p4|b4_p4|b5_p4|b6_p4|b7_p4 \$4042 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1361 \$5127 \$5010 \$5255 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1362 \$5255 \$5011 \$5261 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1363 \$5128 \$5010 \$5259 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1364 \$5259 \$5011 \$4827 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1365 \$3116 \$4145 \$4041 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1366 \$3116 \$4146 \$4041 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1367 \$4541 \$4147 \$3116 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1368 \$4042 \$3612 \$4541 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1369 \$4542 \$3612 \$4041 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1370 \$3328 \$4147 \$4542 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1371 \$4042 \$4145 \$3328 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1372 \$4042 \$4146 \$3328 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1373 b0_r4_b_not \$4145 \$3179 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1374 b0_r4_b_not \$4146 \$3179 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1375 \$4543 \$4147 b0_r4_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1376 \$3178 \$3612 \$4543 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1377 \$4544 \$3612 \$3179 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1378 b0_r4_b \$4147 \$4544 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1379 \$3178 \$4146 b0_r4_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1380 \$3178 \$4145 b0_r4_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1381 \$5072 \$5012 \$4827 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1382 \$5128 \$5013 \$5072 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1383 \$4827 \$5013 \$5073 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1384 \$5074 \$5073 \$5261 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1385 \$5127 \$5072 \$5074 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1386 \$5261 \$5072 \$5075 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1387 \$4046 a3|b0_p3|b1_p3|b2_p3|b3_p3|b5_p3|b6_p3|b7_p3 b2_c2_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1388 b2_c2 a3|b0_p3|b1_p3|b2_p3|b3_p3|b5_p3|b6_p3|b7_p3 \$4047 vdd pfet_03v3
+ L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1389 \$5129 \$5015 \$4151 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1390 \$4151 \$5016 \$5272 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1391 \$5130 \$5015 \$5270 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1392 \$5270 \$5016 \$4829 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1393 \$3117 \$4153 \$4046 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1394 \$3117 \$4152 \$4046 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1395 \$4547 \$4154 \$3117 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1396 \$4047 \$3616 \$4547 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1397 \$4548 \$3616 \$4046 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1398 \$3335 \$4154 \$4548 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1399 \$4047 \$4152 \$3335 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1400 \$4047 \$4153 \$3335 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1401 b2_r3_b_not \$4153 \$3186 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1402 b2_r3_b_not \$4152 \$3186 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1403 \$4549 \$4154 b2_r3_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1404 \$3185 \$3616 \$4549 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1405 \$4550 \$3616 \$3186 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1406 b2_r3_b \$4154 \$4550 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1407 \$3185 \$4153 b2_r3_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1408 \$3185 \$4152 b2_r3_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1409 \$5076 b2_r2_b_not \$4829 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1410 \$5130 b2_r2_b \$5076 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1411 \$4829 b2_r2_b \$5077 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1412 \$5078 \$5077 \$5272 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1413 \$5129 \$5076 \$5078 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1414 \$5272 \$5076 \$5079 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1415 \$4051 a3|b0_p3|b1_p3|b2_p3|b3_p3|b5_p3|b6_p3|b7_p3 b3_c2_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1416 b3_c2 a3|b0_p3|b1_p3|b2_p3|b3_p3|b5_p3|b6_p3|b7_p3 \$4052 vdd pfet_03v3
+ L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1417 \$5080 \$5020 \$4158 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1418 \$4157 \$5021 \$5080 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1419 \$5081 \$5020 \$4157 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1420 \$4158 \$5021 \$5081 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1421 \$5082 \$5020 \$5278 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1422 \$5279 \$5021 \$5082 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1423 \$4831 \$5020 \$5279 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1424 \$5278 \$5021 \$4831 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1425 \$3118 \$4088 \$4051 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1426 \$4052 \$4088 \$3342 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1427 b3_r3_b_not \$4088 \$3120 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1428 \$3119 \$4088 b3_r3_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1429 \$5083 b3_r2_b_not \$4831 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1430 \$5082 b3_r2_b \$5083 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1431 \$5084 b3_r2_b_not \$5082 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1432 \$4831 b3_r2_b \$5084 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1433 \$5085 \$5084 \$5081 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1434 \$5080 \$5083 \$5085 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1435 \$5086 \$5084 \$5080 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1436 \$5081 \$5083 \$5086 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1437 \$4056 b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b4|b4_q7 b4_c2_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1438 \$4056 a3|b0_p3|b1_p3|b2_p3|b3_p3|b5_p3|b6_p3|b7_p3 b4_c2_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1439 \$4557
+ b2_q0_not|b2_q1_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b4_not|b4_q7_not
+ \$4056 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1440 b4_c2
+ a3_not|b0_p3_not|b1_p3_not|b2_p3_not|b3_p3_not|b5_p3_not|b6_p3_not|b7_p3_not
+ \$4557 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1441 \$4558
+ a3_not|b0_p3_not|b1_p3_not|b2_p3_not|b3_p3_not|b5_p3_not|b6_p3_not|b7_p3_not
+ b4_c2_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1442 \$4057
+ b2_q0_not|b2_q1_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b4_not|b4_q7_not
+ \$4558 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1443 b4_c2 a3|b0_p3|b1_p3|b2_p3|b3_p3|b5_p3|b6_p3|b7_p3 \$4057 vdd pfet_03v3
+ L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1444 b4_c2 b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b4|b4_q7 \$4057 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1445 \$5134 \$5025 \$4093 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1446 \$4092 \$5026 \$5134 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1447 \$4093 \$5026 \$5087 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1448 \$5135 \$5025 \$5289 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1449 \$5290 \$5026 \$5135 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1450 \$5289 \$5026 \$4835 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1451 \$3123 \$4095 \$4056 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1452 \$4057 \$4095 \$3349 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1453 b4_r3_b_not \$4094 \$3124 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1454 b4_r3_b_not \$4095 \$3124 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1455 \$4561 \$4160 b4_r3_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1456 \$3195 \$3622 \$4561 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1457 \$4562 \$3622 \$3124 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1458 b4_r3_b \$4160 \$4562 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1459 \$3195 \$4095 b4_r3_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1460 \$3195 \$4094 b4_r3_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1461 \$5088 b4_r2_b_not \$4835 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1462 \$5135 b4_r2_b \$5088 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1463 \$4835 b4_r2_b \$5089 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1464 \$5090 \$5089 \$5087 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1465 \$5134 \$5088 \$5090 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1466 \$5087 \$5088 \$5091 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1467 \$4061 b5|b5_q0|b5_q1|b5_q2|b5_q3|b5_q4|b5_q5|b5_q6|b5_q7 b5_c2_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1468 \$4061 a3|b0_p3|b1_p3|b2_p3|b3_p3|b5_p3|b6_p3|b7_p3 b5_c2_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1469 \$4563
+ b5_not|b5_q0_not|b5_q1_not|b5_q2_not|b5_q3_not|b5_q4_not|b5_q5_not|b5_q6_not|b5_q7_not
+ \$4061 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1470 b5_c2
+ a3_not|b0_p3_not|b1_p3_not|b2_p3_not|b3_p3_not|b5_p3_not|b6_p3_not|b7_p3_not
+ \$4563 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1471 \$4564
+ a3_not|b0_p3_not|b1_p3_not|b2_p3_not|b3_p3_not|b5_p3_not|b6_p3_not|b7_p3_not
+ b5_c2_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1472 \$4062
+ b5_not|b5_q0_not|b5_q1_not|b5_q2_not|b5_q3_not|b5_q4_not|b5_q5_not|b5_q6_not|b5_q7_not
+ \$4564 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1473 b5_c2 b5|b5_q0|b5_q1|b5_q2|b5_q3|b5_q4|b5_q5|b5_q6|b5_q7 \$4062 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1474 b5_c2 a3|b0_p3|b1_p3|b2_p3|b3_p3|b5_p3|b6_p3|b7_p3 \$4062 vdd pfet_03v3
+ L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1475 \$5136 \$5030 \$4164 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1476 \$4163 \$5031 \$5136 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1477 \$4164 \$5031 \$5092 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1478 \$5137 \$5030 \$5299 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1479 \$5300 \$5031 \$5137 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1480 \$5299 \$5031 \$4837 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1481 \$3126 \$4098 \$4061 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1482 \$4062 \$4098 \$3356 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1483 b5_r3_b_not \$4097 \$3127 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1484 b5_r3_b_not \$4098 \$3127 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1485 \$4567 \$4165 b5_r3_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1486 \$3200 \$3624 \$4567 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1487 \$4568 \$3624 \$3127 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1488 b5_r3_b \$4165 \$4568 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1489 \$3200 \$4097 b5_r3_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1490 \$3200 \$4098 b5_r3_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1491 \$5093 b5_r2_b_not \$4837 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1492 \$5137 b5_r2_b \$5093 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1493 \$4837 b5_r2_b \$5094 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1494 \$5095 \$5094 \$5092 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1495 \$5136 \$5093 \$5095 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1496 \$5092 \$5093 \$5096 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1497 \$4066 a3|b0_p3|b1_p3|b2_p3|b3_p3|b5_p3|b6_p3|b7_p3 b6_c2_not|b6_c3_not
+ vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1498 b6_c2|b6_c3 a3|b0_p3|b1_p3|b2_p3|b3_p3|b5_p3|b6_p3|b7_p3 \$4067 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1499 \$5138 \$5035 \$4169 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1500 \$4168 \$5036 \$5138 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1501 \$4169 \$5036 \$5097 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1502 \$5139 \$5035 \$5308 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1503 \$5309 \$5036 \$5139 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1504 \$5308 \$5036 \$4839 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1505 \$3129 \$4101 \$4066 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1506 \$4067 \$4101 \$3364 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1507 b6_r3_b_not \$4101 \$3130 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1508 b6_r3_b_not \$4100 \$3130 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1509 \$4573 \$4170 b6_r3_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1510 \$3205 \$3626 \$4573 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1511 \$4574 \$3626 \$3130 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1512 b6_r3_b \$4170 \$4574 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1513 \$3205 \$4101 b6_r3_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1514 \$3205 \$4100 b6_r3_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1515 \$5098 b6_r2_b_not \$4839 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1516 \$5139 b6_r2_b \$5098 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1517 \$4839 b6_r2_b \$5099 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1518 \$5100 \$5099 \$5097 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1519 \$5138 \$5098 \$5100 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1520 \$5097 \$5098 \$5101 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1521 \$4071 a3|b0_p3|b1_p3|b2_p3|b3_p3|b5_p3|b6_p3|b7_p3 b6_c2_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1522 b6_c2 a3|b0_p3|b1_p3|b2_p3|b3_p3|b5_p3|b6_p3|b7_p3 \$4072 vdd pfet_03v3
+ L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1523 \$5140 \$5040 \$4174 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1524 \$4173 \$5041 \$5140 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1525 \$4174 \$5041 \$5102 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1526 \$5141 \$5040 \$5318 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1527 \$5319 \$5041 \$5141 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1528 \$5318 \$5041 \$4841 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1529 \$3132 \$4104 \$4071 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1530 \$4072 \$4104 \$3371 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1531 \$4073 \$4103 \$3133 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1532 \$4073 \$4104 \$3133 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1533 \$4579 \$4175 \$4073 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1534 \$3210 \$3628 \$4579 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1535 \$4580 \$3628 \$3133 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1536 \$4074 \$4175 \$4580 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1537 \$3210 \$4103 \$4074 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1538 \$3210 \$4104 \$4074 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1539 \$5103 \$5042 \$4841 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1540 \$5141 \$5043 \$5103 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1541 \$4841 \$5043 \$5104 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1542 p9 \$5104 \$5102 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$1543 \$5140 \$5103 p9 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$1544 \$5102 \$5103 p9_not vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1545 \$5255 b1|b1_q0|b1_q1|b1_q2|b1_q3|b1_q4|b1_q5|b1_q6|b1_q7 b1_c2_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1546 \$5508
+ b1_not|b1_q0_not|b1_q1_not|b1_q2_not|b1_q3_not|b1_q4_not|b1_q5_not|b1_q6_not|b1_q7_not
+ \$5255 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1547 b1_c2
+ a2_not|b0_p2_not|b1_p2_not|b2_p2_not|b3_p2_not|b5_p2_not|b6_p2_not|b7_p2_not
+ \$5508 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1548 \$5509
+ a2_not|b0_p2_not|b1_p2_not|b2_p2_not|b3_p2_not|b5_p2_not|b6_p2_not|b7_p2_not
+ b1_c2_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1549 \$5008
+ b1_not|b1_q0_not|b1_q1_not|b1_q2_not|b1_q3_not|b1_q4_not|b1_q5_not|b1_q6_not|b1_q7_not
+ \$5509 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1550 b1_c2 b1|b1_q0|b1_q1|b1_q2|b1_q3|b1_q4|b1_q5|b1_q6|b1_q7 \$5008 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1551 \$5010 b0|b0_q0|b0_q1|b0_q2|b0_q3|b0_q4|b0_q5|b0_q6|b0_q7 b0_c3_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1552 \$5510
+ b0_not|b0_q0_not|b0_q1_not|b0_q3_not|b0_q4_not|b0_q5_not|b0_q6_not|b0_q7_not|b1_q2_not
+ \$5010 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1553 b0_c3
+ a3_not|b0_p3_not|b1_p3_not|b2_p3_not|b3_p3_not|b5_p3_not|b6_p3_not|b7_p3_not
+ \$5510 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1554 \$5511
+ a3_not|b0_p3_not|b1_p3_not|b2_p3_not|b3_p3_not|b5_p3_not|b6_p3_not|b7_p3_not
+ b0_c3_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1555 \$5011
+ b0_not|b0_q0_not|b0_q1_not|b0_q3_not|b0_q4_not|b0_q5_not|b0_q6_not|b0_q7_not|b1_q2_not
+ \$5511 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1556 b0_c3 b0|b0_q0|b0_q1|b0_q2|b0_q3|b0_q4|b0_q5|b0_q6|b0_q7 \$5011 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1557 \$5008 \$5011 \$5127 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1558 \$5261 \$5010 \$5008 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1559 \$5260 \$5011 \$5128 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1560 \$4827 \$5010 \$5260 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1561 \$5073 \$5012 \$5128 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1562 \$5075 \$5073 \$5127 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1563 \$5015 b2|b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7 b2_c2_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1564 \$5516
+ b2_not|b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not
+ \$5015 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1565 b2_c2
+ a2_not|b0_p2_not|b1_p2_not|b2_p2_not|b3_p2_not|b5_p2_not|b6_p2_not|b7_p2_not
+ \$5516 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1566 \$5517
+ a2_not|b0_p2_not|b1_p2_not|b2_p2_not|b3_p2_not|b5_p2_not|b6_p2_not|b7_p2_not
+ b2_c2_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1567 \$5016
+ b2_not|b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not
+ \$5517 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1568 b2_c2 b2|b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7 \$5016 vdd pfet_03v3
+ L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1569 \$4150 \$5016 \$5129 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1570 \$5272 \$5015 \$4150 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1571 \$5271 \$5016 \$5130 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1572 \$4829 \$5015 \$5271 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1573 \$5077 b2_r2_b_not \$5130 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1574 \$5079 \$5077 \$5129 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1575 \$5020
+ b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b3|b3_q0|b3_q1|b3_q2|b3_q3|b3_q4|b3_q5|b3_q6|b3_q7
+ b3_c2_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1576 \$5522
+ b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b3_not|b3_q0_not|b3_q1_not|b3_q2_not|b3_q3_not|b3_q4_not|b3_q5_not|b3_q6_not|b3_q7_not
+ \$5020 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1577 b3_c2
+ a2_not|b0_p2_not|b1_p2_not|b2_p2_not|b3_p2_not|b5_p2_not|b6_p2_not|b7_p2_not
+ \$5522 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1578 \$5523
+ a2_not|b0_p2_not|b1_p2_not|b2_p2_not|b3_p2_not|b5_p2_not|b6_p2_not|b7_p2_not
+ b3_c2_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1579 \$5021
+ b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b3_not|b3_q0_not|b3_q1_not|b3_q2_not|b3_q3_not|b3_q4_not|b3_q5_not|b3_q6_not|b3_q7_not
+ \$5523 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1580 b3_c2
+ b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b3|b3_q0|b3_q1|b3_q2|b3_q3|b3_q4|b3_q5|b3_q6|b3_q7
+ \$5021 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1581 \$4089 \$5080 \$5020 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1582 \$5524 \$5081 \$4089 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1583 \$5021 \$4831 \$5524 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1584 \$5525 \$4831 \$5020 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1585 \$4309 \$5081 \$5525 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1586 \$5021 \$5080 \$4309 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1587 b3_r2_b_not \$5080 \$4091 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1588 \$5526 \$5081 b3_r2_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1589 \$4090 \$4831 \$5526 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1590 \$5527 \$4831 \$4091 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1591 b3_r2_b \$5081 \$5527 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1592 \$4090 \$5080 b3_r2_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1593 \$5025 b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b4|b4_q7 b4_c2_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1594 \$5528
+ b2_q0_not|b2_q1_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b4_not|b4_q7_not
+ \$5025 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1595 b4_c2
+ a2_not|b0_p2_not|b1_p2_not|b2_p2_not|b3_p2_not|b5_p2_not|b6_p2_not|b7_p2_not
+ \$5528 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1596 \$5529
+ a2_not|b0_p2_not|b1_p2_not|b2_p2_not|b3_p2_not|b5_p2_not|b6_p2_not|b7_p2_not
+ b4_c2_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1597 \$5026
+ b2_q0_not|b2_q1_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b4_not|b4_q7_not
+ \$5529 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1598 b4_c2 b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b4|b4_q7 \$5026 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1599 \$5087 \$5025 \$4092 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1600 \$4835 \$5025 \$5290 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1601 \$5089 b4_r2_b_not \$5135 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1602 \$5091 \$5089 \$5134 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1603 \$5030 b5|b5_q0|b5_q1|b5_q2|b5_q3|b5_q4|b5_q5|b5_q6|b5_q7 b5_c2_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1604 \$5534
+ b5_not|b5_q0_not|b5_q1_not|b5_q2_not|b5_q3_not|b5_q4_not|b5_q5_not|b5_q6_not|b5_q7_not
+ \$5030 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1605 b5_c2
+ a2_not|b0_p2_not|b1_p2_not|b2_p2_not|b3_p2_not|b5_p2_not|b6_p2_not|b7_p2_not
+ \$5534 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1606 \$5535
+ a2_not|b0_p2_not|b1_p2_not|b2_p2_not|b3_p2_not|b5_p2_not|b6_p2_not|b7_p2_not
+ b5_c2_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1607 \$5031
+ b5_not|b5_q0_not|b5_q1_not|b5_q2_not|b5_q3_not|b5_q4_not|b5_q5_not|b5_q6_not|b5_q7_not
+ \$5535 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1608 b5_c2 b5|b5_q0|b5_q1|b5_q2|b5_q3|b5_q4|b5_q5|b5_q6|b5_q7 \$5031 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1609 \$5092 \$5030 \$4163 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1610 \$4837 \$5030 \$5300 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1611 \$5094 b5_r2_b_not \$5137 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1612 \$5096 \$5094 \$5136 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1613 \$5035 b6|b6_q0|b6_q1|b6_q2|b6_q3|b6_q4|b6_q5|b6_q6|b6_q7 b6_c2_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1614 \$5540
+ b6_not|b6_q0_not|b6_q1_not|b6_q2_not|b6_q3_not|b6_q4_not|b6_q5_not|b6_q6_not|b6_q7_not
+ \$5035 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1615 b6_c2
+ a2_not|b0_p2_not|b1_p2_not|b2_p2_not|b3_p2_not|b5_p2_not|b6_p2_not|b7_p2_not
+ \$5540 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1616 \$5541
+ a2_not|b0_p2_not|b1_p2_not|b2_p2_not|b3_p2_not|b5_p2_not|b6_p2_not|b7_p2_not
+ b6_c2_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1617 \$5036
+ b6_not|b6_q0_not|b6_q1_not|b6_q2_not|b6_q3_not|b6_q4_not|b6_q5_not|b6_q6_not|b6_q7_not
+ \$5541 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1618 b6_c2 b6|b6_q0|b6_q1|b6_q2|b6_q3|b6_q4|b6_q5|b6_q6|b6_q7 \$5036 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1619 \$5097 \$5035 \$4168 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1620 \$4839 \$5035 \$5309 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1621 \$5099 b6_r2_b_not \$5139 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1622 \$5101 \$5099 \$5138 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1623 \$5040 b1_q3|b7|b7_q0|b7_q1|b7_q2|b7_q4|b7_q5|b7_q6|b7_q7 b6_c2_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1624 \$5546
+ b7_not|b7_q0_not|b7_q1_not|b7_q2_not|b7_q3_not|b7_q4_not|b7_q5_not|b7_q6_not|b7_q7_not
+ \$5040 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1625 b6_c2
+ a2_not|b0_p2_not|b1_p2_not|b2_p2_not|b3_p2_not|b5_p2_not|b6_p2_not|b7_p2_not
+ \$5546 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1626 \$5547
+ a2_not|b0_p2_not|b1_p2_not|b2_p2_not|b3_p2_not|b5_p2_not|b6_p2_not|b7_p2_not
+ b6_c2_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1627 \$5041
+ b7_not|b7_q0_not|b7_q1_not|b7_q2_not|b7_q3_not|b7_q4_not|b7_q5_not|b7_q6_not|b7_q7_not
+ \$5547 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1628 b6_c2 b1_q3|b7|b7_q0|b7_q1|b7_q2|b7_q4|b7_q5|b7_q6|b7_q7 \$5041 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1629 \$5102 \$5040 \$4173 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1630 \$4841 \$5040 \$5319 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1631 \$5104 \$5042 \$5141 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1632 p9_not \$5104 \$5140 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1633 \$5255 a2|b0_p2|b1_p2|b2_p2|b3_p2|b4_p2|b5_p2|b6_p2|b7_p2 b1_c2_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1634 b1_c2 a2|b0_p2|b1_p2|b2_p2|b3_p2|b4_p2|b5_p2|b6_p2|b7_p2 \$5008 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1635 \$5010 a3|b0_p3|b1_p3|b2_p3|b3_p3|b5_p3|b6_p3|b7_p3 b0_c3_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1636 b0_c3 a3|b0_p3|b1_p3|b2_p3|b3_p3|b5_p3|b6_p3|b7_p3 \$5011 vdd pfet_03v3
+ L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1637 \$4085 \$5127 \$5010 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1638 \$4085 \$5128 \$5010 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1639 \$5512 \$5261 \$4085 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1640 \$5011 \$4827 \$5512 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1641 \$5513 \$4827 \$5010 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1642 \$4293 \$5261 \$5513 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1643 \$5011 \$5128 \$4293 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1644 \$5011 \$5127 \$4293 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1645 \$5012 \$5127 \$4149 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1646 \$5012 \$5128 \$4149 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1647 \$5514 \$5261 \$5012 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1648 \$4148 \$4827 \$5514 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1649 \$5515 \$4827 \$4149 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1650 \$5013 \$5261 \$5515 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1651 \$4148 \$5128 \$5013 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1652 \$4148 \$5127 \$5013 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1653 \$6062 \$5950 \$5798 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1654 \$6061 \$5951 \$6062 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1655 \$5798 \$5951 \$6063 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1656 \$6064 \$6063 \$6060 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1657 \$6059 \$6062 \$6064 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1658 \$6060 \$6062 \$6065 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1659 \$5015 a2|b0_p2|b1_p2|b2_p2|b3_p2|b4_p2|b5_p2|b6_p2|b7_p2 b2_c2_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1660 b2_c2 a2|b0_p2|b1_p2|b2_p2|b3_p2|b4_p2|b5_p2|b6_p2|b7_p2 \$5016 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1661 \$4086 \$5130 \$5015 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1662 \$4086 \$5129 \$5015 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1663 \$5518 \$5272 \$4086 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1664 \$5016 \$4829 \$5518 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1665 \$5519 \$4829 \$5015 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1666 \$4301 \$5272 \$5519 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1667 \$5016 \$5129 \$4301 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1668 \$5016 \$5130 \$4301 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1669 b2_r2_b_not \$5130 \$4156 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1670 b2_r2_b_not \$5129 \$4156 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1671 \$5520 \$5272 b2_r2_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1672 \$4155 \$4829 \$5520 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1673 \$5521 \$4829 \$4156 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1674 b2_r2_b \$5272 \$5521 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1675 \$4155 \$5129 b2_r2_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1676 \$4155 \$5130 b2_r2_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1677 \$6069 b2_r1_b_not \$5800 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1678 \$6068 b2_r1_b \$6069 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1679 \$5800 b2_r1_b \$6070 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1680 \$6071 \$6070 \$6067 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1681 \$6066 \$6069 \$6071 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1682 \$6067 \$6069 \$6072 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1683 \$5020 a2|b0_p2|b1_p2|b2_p2|b3_p2|b4_p2|b5_p2|b6_p2|b7_p2 b3_c2_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1684 b3_c2 a2|b0_p2|b1_p2|b2_p2|b3_p2|b4_p2|b5_p2|b6_p2|b7_p2 \$5021 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1685 \$6073 \$5956 \$5079 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1686 \$5079 \$6000 \$6074 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1687 \$6075 \$5956 \$6180 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1688 \$6180 \$6000 \$5802 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1689 \$4089 \$5082 \$5020 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1690 \$5021 \$5082 \$4309 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1691 b3_r2_b_not \$5082 \$4091 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1692 \$4090 \$5082 b3_r2_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1693 \$6076 b3_r1_b_not \$5802 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1694 \$6075 b3_r1_b \$6076 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1695 \$6077 b3_r1_b_not \$6075 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1696 \$5802 b3_r1_b \$6077 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1697 \$6078 \$6077 \$6074 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1698 \$6073 \$6076 \$6078 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1699 \$6079 \$6077 \$6073 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1700 \$6074 \$6076 \$6079 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1701 \$5025 a2|b0_p2|b1_p2|b2_p2|b3_p2|b4_p2|b5_p2|b6_p2|b7_p2 b4_c2_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1702 b4_c2 a2|b0_p2|b1_p2|b2_p2|b3_p2|b4_p2|b5_p2|b6_p2|b7_p2 \$5026 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1703 \$4096 \$5134 \$5025 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1704 \$4096 \$5135 \$5025 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1705 \$5530 \$5087 \$4096 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1706 \$5026 \$4835 \$5530 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1707 \$5531 \$4835 \$5025 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1708 \$4317 \$5087 \$5531 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1709 \$5026 \$5134 \$4317 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1710 \$5026 \$5135 \$4317 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1711 b4_r2_b_not \$5134 \$4162 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1712 b4_r2_b_not \$5135 \$4162 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1713 \$5532 \$5087 b4_r2_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1714 \$4161 \$4835 \$5532 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1715 \$5533 \$4835 \$4162 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1716 b4_r2_b \$5087 \$5533 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1717 \$4161 \$5135 b4_r2_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1718 \$4161 \$5134 b4_r2_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1719 \$6083 b4_r1_b_not \$5804 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1720 \$6082 b4_r1_b \$6083 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1721 \$6084 b4_r1_b_not \$6082 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1722 \$5804 b4_r1_b \$6084 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1723 \$6085 \$6084 \$6081 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1724 \$6080 \$6083 \$6085 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1725 \$6086 \$6084 \$6080 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1726 \$6081 \$6083 \$6086 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1727 \$5030 a2|b0_p2|b1_p2|b2_p2|b3_p2|b4_p2|b5_p2|b6_p2|b7_p2 b5_c2_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1728 b5_c2 a2|b0_p2|b1_p2|b2_p2|b3_p2|b4_p2|b5_p2|b6_p2|b7_p2 \$5031 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1729 \$4099 \$5136 \$5030 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1730 \$4099 \$5137 \$5030 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1731 \$5536 \$5092 \$4099 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1732 \$5031 \$4837 \$5536 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1733 \$5537 \$4837 \$5030 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1734 \$4325 \$5092 \$5537 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1735 \$5031 \$5136 \$4325 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1736 \$5031 \$5137 \$4325 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1737 b5_r2_b_not \$5137 \$4167 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1738 b5_r2_b_not \$5136 \$4167 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1739 \$5538 \$5092 b5_r2_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1740 \$4166 \$4837 \$5538 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1741 \$5539 \$4837 \$4167 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1742 b5_r2_b \$5092 \$5539 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1743 \$4166 \$5136 b5_r2_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1744 \$4166 \$5137 b5_r2_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1745 \$6090 b5_r1_b_not \$5806 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1746 \$6089 b5_r1_b \$6090 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1747 \$6091 b5_r1_b_not \$6089 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1748 \$5806 b5_r1_b \$6091 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1749 \$6092 \$6091 \$6088 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1750 \$6087 \$6090 \$6092 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1751 \$6093 \$6091 \$6087 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1752 \$6088 \$6090 \$6093 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1753 \$5035 a2|b0_p2|b1_p2|b2_p2|b3_p2|b4_p2|b5_p2|b6_p2|b7_p2 b6_c2_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1754 b6_c2 a2|b0_p2|b1_p2|b2_p2|b3_p2|b4_p2|b5_p2|b6_p2|b7_p2 \$5036 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1755 \$4102 \$5139 \$5035 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1756 \$4102 \$5138 \$5035 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1757 \$5542 \$5097 \$4102 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1758 \$5036 \$4839 \$5542 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1759 \$5543 \$4839 \$5035 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1760 \$4332 \$5097 \$5543 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1761 \$5036 \$5139 \$4332 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1762 \$5036 \$5138 \$4332 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1763 b6_r2_b_not \$5139 \$4172 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1764 b6_r2_b_not \$5138 \$4172 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1765 \$5544 \$5097 b6_r2_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1766 \$4171 \$4839 \$5544 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1767 \$5545 \$4839 \$4172 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1768 b6_r2_b \$5097 \$5545 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1769 \$4171 \$5138 b6_r2_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1770 \$4171 \$5139 b6_r2_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1771 \$6097 b6_r1_b_not \$5808 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1772 \$6096 b6_r1_b \$6097 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1773 \$6098 b6_r1_b_not \$6096 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1774 \$5808 b6_r1_b \$6098 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1775 \$6099 \$6098 \$6095 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1776 \$6094 \$6097 \$6099 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1777 \$6100 \$6098 \$6094 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1778 \$6095 \$6097 \$6100 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1779 \$5040 a2|b0_p2|b1_p2|b2_p2|b3_p2|b4_p2|b5_p2|b6_p2|b7_p2 b6_c2_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1780 b6_c2 a2|b0_p2|b1_p2|b2_p2|b3_p2|b4_p2|b5_p2|b6_p2|b7_p2 \$5041 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1781 \$4105 \$5140 \$5040 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1782 \$4105 \$5141 \$5040 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1783 \$5548 \$5102 \$4105 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1784 \$5041 \$4841 \$5548 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1785 \$5549 \$4841 \$5040 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1786 \$4340 \$5102 \$5549 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1787 \$5041 \$5140 \$4340 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1788 \$5041 \$5141 \$4340 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1789 \$5042 \$5141 \$4177 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1790 \$5042 \$5140 \$4177 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1791 \$5550 \$5102 \$5042 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1792 \$4176 \$4841 \$5550 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1793 \$5551 \$4841 \$4177 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1794 \$5043 \$5102 \$5551 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1795 \$4176 \$5141 \$5043 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1796 \$4176 \$5140 \$5043 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1797 \$6104 \$5970 \$5810 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1798 \$6103 \$5971 \$6104 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1799 \$6105 \$5970 \$6103 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1800 \$5810 \$5971 \$6105 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1801 p8 \$6105 \$6102 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$1802 \$6101 \$6104 p8 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$1803 p8_not \$6105 \$6101 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1804 \$6102 \$6104 p8_not vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1805 \$6059 \$5995 \$6409 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1806 \$5948 \$5996 \$6059 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1807 \$6060 \$5995 \$5948 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1808 \$6409 \$5996 \$6060 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1809 \$6061 \$5995 \$6164 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1810 \$6411 \$5996 \$6061 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1811 \$5798 \$5995 \$6411 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1812 \$6164 \$5996 \$5798 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1813 \$6063 \$5950 \$6061 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1814 \$6065 \$6063 \$6059 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1815 \$6066 \$5998 \$5075 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1816 \$5074 \$5999 \$6066 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1817 \$6067 \$5998 \$5074 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1818 \$5075 \$5999 \$6067 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1819 \$6068 \$5998 \$6172 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1820 \$6413 \$5999 \$6068 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1821 \$5800 \$5998 \$6413 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1822 \$6172 \$5999 \$5800 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1823 \$6070 b2_r1_b_not \$6068 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1824 \$6072 \$6070 \$6066 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1825 \$5078 \$6000 \$6073 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1826 \$6074 \$5956 \$5078 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1827 \$6416 \$6000 \$6075 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1828 \$5802 \$5956 \$6416 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1829 \$6080 \$6002 \$5086 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1830 \$5085 \$6003 \$6080 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1831 \$6081 \$6002 \$5085 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1832 \$5086 \$6003 \$6081 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1833 \$6082 \$6002 \$6188 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1834 \$6419 \$6003 \$6082 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1835 \$5804 \$6002 \$6419 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1836 \$6188 \$6003 \$5804 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1837 \$6087 \$6005 \$5091 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1838 \$5090 \$6006 \$6087 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1839 \$6088 \$6005 \$5090 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1840 \$5091 \$6006 \$6088 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1841 \$6089 \$6005 \$6196 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1842 \$6422 \$6006 \$6089 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1843 \$5806 \$6005 \$6422 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1844 \$6196 \$6006 \$5806 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1845 \$6094 \$6008 \$5096 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1846 \$5095 \$6009 \$6094 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1847 \$6095 \$6008 \$5095 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1848 \$5096 \$6009 \$6095 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1849 \$6096 \$6008 \$6203 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1850 \$6425 \$6009 \$6096 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1851 \$5808 \$6008 \$6425 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1852 \$6203 \$6009 \$5808 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1853 \$6101 \$6011 \$5101 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1854 \$5100 \$6012 \$6101 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1855 \$6102 \$6011 \$5100 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1856 \$5101 \$6012 \$6102 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1857 \$6103 \$6011 \$6211 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1858 \$6427 \$6012 \$6103 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1859 \$5810 \$6011 \$6427 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1860 \$6211 \$6012 \$5810 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1861 \$6409 b1|b1_q0|b1_q1|b1_q2|b1_q3|b1_q4|b1_q5|b1_q6|b1_q7 b1_c1_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1862 \$6476
+ b1_not|b1_q0_not|b1_q1_not|b1_q2_not|b1_q3_not|b1_q4_not|b1_q5_not|b1_q6_not|b1_q7_not
+ \$6409 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1863 b1_c1
+ a1_not|b0_p1_not|b1_p1_not|b2_p1_not|b3_p1_not|b4_p1_not|b5_p1_not|b6_p1_not|b7_p1_not
+ \$6476 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1864 \$6477
+ a1_not|b0_p1_not|b1_p1_not|b2_p1_not|b3_p1_not|b4_p1_not|b5_p1_not|b6_p1_not|b7_p1_not
+ b1_c1_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1865 \$5948
+ b1_not|b1_q0_not|b1_q1_not|b1_q2_not|b1_q3_not|b1_q4_not|b1_q5_not|b1_q6_not|b1_q7_not
+ \$6477 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1866 b1_c1 b1|b1_q0|b1_q1|b1_q2|b1_q3|b1_q4|b1_q5|b1_q6|b1_q7 \$5948 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1867 \$5995 b0|b0_q0|b0_q1|b0_q2|b0_q3|b0_q4|b0_q5|b0_q6|b0_q7 b0_c2_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1868 \$6492
+ b0_not|b0_q0_not|b0_q1_not|b0_q3_not|b0_q4_not|b0_q5_not|b0_q6_not|b0_q7_not|b1_q2_not
+ \$5995 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1869 b0_c2
+ a2_not|b0_p2_not|b1_p2_not|b2_p2_not|b3_p2_not|b5_p2_not|b6_p2_not|b7_p2_not
+ \$6492 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1870 \$6493
+ a2_not|b0_p2_not|b1_p2_not|b2_p2_not|b3_p2_not|b5_p2_not|b6_p2_not|b7_p2_not
+ b0_c2_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1871 \$5996
+ b0_not|b0_q0_not|b0_q1_not|b0_q3_not|b0_q4_not|b0_q5_not|b0_q6_not|b0_q7_not|b1_q2_not
+ \$6493 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1872 b0_c2 b0|b0_q0|b0_q1|b0_q2|b0_q3|b0_q4|b0_q5|b0_q6|b0_q7 \$5996 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1873 \$5259 \$6059 \$5995 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1874 \$6494 \$6060 \$5259 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1875 \$5996 \$5798 \$6494 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1876 \$6495 \$5798 \$5995 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1877 \$5260 \$6060 \$6495 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1878 \$5996 \$6059 \$5260 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1879 \$5950 \$6059 \$5073 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1880 \$6478 \$6060 \$5950 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1881 \$5072 \$5798 \$6478 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1882 \$6479 \$5798 \$5073 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1883 \$5951 \$6060 \$6479 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1884 \$5072 \$6059 \$5951 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1885 \$5998 b2|b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7 b2_c1_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1886 \$6496
+ b2_not|b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not
+ \$5998 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1887 b2_c1
+ a1_not|b0_p1_not|b1_p1_not|b2_p1_not|b3_p1_not|b4_p1_not|b5_p1_not|b6_p1_not|b7_p1_not
+ \$6496 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1888 \$6497
+ a1_not|b0_p1_not|b1_p1_not|b2_p1_not|b3_p1_not|b4_p1_not|b5_p1_not|b6_p1_not|b7_p1_not
+ b2_c1_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1889 \$5999
+ b2_not|b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not
+ \$6497 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1890 b2_c1 b2|b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7 \$5999 vdd pfet_03v3
+ L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1891 \$5270 \$6066 \$5998 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1892 \$6498 \$6067 \$5270 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1893 \$5999 \$5800 \$6498 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1894 \$6499 \$5800 \$5998 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1895 \$5271 \$6067 \$6499 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1896 \$5999 \$6066 \$5271 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1897 b2_r1_b_not \$6066 \$5077 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1898 \$6480 \$6067 b2_r1_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1899 \$5076 \$5800 \$6480 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1900 \$6481 \$5800 \$5077 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1901 b2_r1_b \$6067 \$6481 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1902 \$5076 \$6066 b2_r1_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1903 \$5956
+ b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b3|b3_q0|b3_q1|b3_q2|b3_q3|b3_q4|b3_q5|b3_q6|b3_q7
+ b2_c1_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1904 \$6500
+ b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b3_not|b3_q0_not|b3_q1_not|b3_q2_not|b3_q3_not|b3_q4_not|b3_q5_not|b3_q6_not|b3_q7_not
+ \$5956 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1905 b3_c1
+ a1_not|b0_p1_not|b1_p1_not|b2_p1_not|b3_p1_not|b4_p1_not|b5_p1_not|b6_p1_not|b7_p1_not
+ \$6500 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1906 \$6501
+ a1_not|b0_p1_not|b1_p1_not|b2_p1_not|b3_p1_not|b4_p1_not|b5_p1_not|b6_p1_not|b7_p1_not
+ b2_c1_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1907 \$6000
+ b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b3_not|b3_q0_not|b3_q1_not|b3_q2_not|b3_q3_not|b3_q4_not|b3_q5_not|b3_q6_not|b3_q7_not
+ \$6501 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1908 b3_c1
+ b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b3|b3_q0|b3_q1|b3_q2|b3_q3|b3_q4|b3_q5|b3_q6|b3_q7
+ \$6000 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1909 \$5278 \$6073 \$5956 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1910 \$6503 \$6074 \$5278 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1911 \$6000 \$5802 \$6503 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1912 \$6504 \$5802 \$5956 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1913 \$5279 \$6074 \$6504 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1914 \$6000 \$6073 \$5279 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1915 b3_r1_b_not \$6073 \$5084 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1916 \$6482 \$6074 b3_r1_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1917 \$5083 \$5802 \$6482 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1918 \$6483 \$5802 \$5084 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1919 b3_r1_b \$6074 \$6483 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1920 \$5083 \$6073 b3_r1_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1921 \$5289 \$6080 \$6002 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1922 \$6508 \$6081 \$5289 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1923 \$6003 \$5804 \$6508 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1924 \$6509 \$5804 \$6002 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1925 \$5290 \$6081 \$6509 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1926 \$6003 \$6080 \$5290 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1927 b4_r1_b_not \$6080 \$5089 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1928 \$6484 \$6081 b4_r1_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1929 \$5088 \$5804 \$6484 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1930 \$6485 \$5804 \$5089 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1931 b4_r1_b \$6081 \$6485 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1932 \$5088 \$6080 b4_r1_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1933 \$5299 \$6087 \$6005 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1934 \$6513 \$6088 \$5299 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1935 \$6006 \$5806 \$6513 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1936 \$6514 \$5806 \$6005 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1937 \$5300 \$6088 \$6514 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1938 \$6006 \$6087 \$5300 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1939 b5_r1_b_not \$6087 \$5094 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1940 \$6486 \$6088 b5_r1_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1941 \$5093 \$5806 \$6486 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1942 \$6487 \$5806 \$5094 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1943 b5_r1_b \$6088 \$6487 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1944 \$5093 \$6087 b5_r1_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1945 \$6008 b6|b6_q0|b6_q1|b6_q2|b6_q3|b6_q4|b6_q5|b6_q6|b6_q7 b6_c1_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1946 \$6515
+ b6_not|b6_q0_not|b6_q1_not|b6_q2_not|b6_q3_not|b6_q4_not|b6_q5_not|b6_q6_not|b6_q7_not
+ \$6008 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1947 b6_c1
+ a1_not|b0_p1_not|b1_p1_not|b2_p1_not|b3_p1_not|b4_p1_not|b5_p1_not|b6_p1_not|b7_p1_not
+ \$6515 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1948 \$6516
+ a1_not|b0_p1_not|b1_p1_not|b2_p1_not|b3_p1_not|b4_p1_not|b5_p1_not|b6_p1_not|b7_p1_not
+ b6_c1_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1949 \$6009
+ b6_not|b6_q0_not|b6_q1_not|b6_q2_not|b6_q3_not|b6_q4_not|b6_q5_not|b6_q6_not|b6_q7_not
+ \$6516 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1950 b6_c1 b6|b6_q0|b6_q1|b6_q2|b6_q3|b6_q4|b6_q5|b6_q6|b6_q7 \$6009 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1951 \$5308 \$6094 \$6008 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1952 \$6518 \$6095 \$5308 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1953 \$6009 \$5808 \$6518 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1954 \$6519 \$5808 \$6008 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1955 \$5309 \$6095 \$6519 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1956 \$6009 \$6094 \$5309 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1957 b6_r1_b_not \$6094 \$5099 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1958 \$6488 \$6095 b6_r1_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$1959 \$5098 \$5808 \$6488 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1960 \$6489 \$5808 \$5099 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1961 b6_r1_b \$6095 \$6489 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1962 \$5098 \$6094 b6_r1_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1963 \$6011 b1_q3|b7|b7_q0|b7_q1|b7_q2|b7_q4|b7_q5|b7_q6|b7_q7 \$6010 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1964 \$6520
+ b7_not|b7_q0_not|b7_q1_not|b7_q2_not|b7_q3_not|b7_q4_not|b7_q5_not|b7_q6_not|b7_q7_not
+ \$6011 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1965 b6_c1
+ a1_not|b0_p1_not|b1_p1_not|b2_p1_not|b3_p1_not|b4_p1_not|b5_p1_not|b6_p1_not|b7_p1_not
+ \$6520 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1966 \$6521
+ a1_not|b0_p1_not|b1_p1_not|b2_p1_not|b3_p1_not|b4_p1_not|b5_p1_not|b6_p1_not|b7_p1_not
+ \$6010 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1967 \$6012
+ b7_not|b7_q0_not|b7_q1_not|b7_q2_not|b7_q3_not|b7_q4_not|b7_q5_not|b7_q6_not|b7_q7_not
+ \$6521 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1968 b6_c1 b1_q3|b7|b7_q0|b7_q1|b7_q2|b7_q4|b7_q5|b7_q6|b7_q7 \$6012 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1969 \$5318 \$6101 \$6011 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1970 \$6523 \$6102 \$5318 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1971 \$6012 \$5810 \$6523 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1972 \$6524 \$5810 \$6011 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1973 \$5319 \$6102 \$6524 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1974 \$6012 \$6101 \$5319 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1975 \$5970 \$6101 \$5104 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1976 \$6490 \$6102 \$5970 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1977 \$5103 \$5810 \$6490 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1978 \$6491 \$5810 \$5104 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1979 \$5971 \$6102 \$6491 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1980 \$5103 \$6101 \$5971 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$1981 \$6409 a1|b0_p1|b1_p1|b2_p1|b3_p1|b4_p1|b5_p1|b6_p1|b7_p1 b1_c1_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1982 \$6929 b1|b1_q0|b1_q1|b1_q2|b1_q3|b1_q4|b1_q5|b1_q6|b1_q7 b1_c0_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1983 \$7445
+ b1_not|b1_q0_not|b1_q1_not|b1_q2_not|b1_q3_not|b1_q4_not|b1_q5_not|b1_q6_not|b1_q7_not
+ \$6929 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1984 b1_c0
+ a0_not|b0_p0_not|b1_p0_not|b2_p0_not|b3_p0_not|b5_p0_not|b6_p0_not|b7_p0_not
+ \$7445 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1985 \$7446
+ a0_not|b0_p0_not|b1_p0_not|b2_p0_not|b3_p0_not|b5_p0_not|b6_p0_not|b7_p0_not
+ b1_c0_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1986 \$6930
+ b1_not|b1_q0_not|b1_q1_not|b1_q2_not|b1_q3_not|b1_q4_not|b1_q5_not|b1_q6_not|b1_q7_not
+ \$7446 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1987 b1_c1 a1|b0_p1|b1_p1|b2_p1|b3_p1|b4_p1|b5_p1|b6_p1|b7_p1 \$5948 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1988 b1_c0 b1|b1_q0|b1_q1|b1_q2|b1_q3|b1_q4|b1_q5|b1_q6|b1_q7 \$6930 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1989 \$5995 a2|b0_p2|b1_p2|b2_p2|b3_p2|b4_p2|b5_p2|b6_p2|b7_p2 b0_c2_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1990 b0_c2 a2|b0_p2|b1_p2|b2_p2|b3_p2|b4_p2|b5_p2|b6_p2|b7_p2 \$5996 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$1991 \$6997 \$7232 \$6929 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1992 \$6930 \$6932 \$6997 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1993 \$6998 \$7232 \$6930 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1994 \$6929 \$6932 \$6998 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1995 \$6999 \$7232 x0_c0_f_not vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$1996 x0_c0_f \$6932 \$6999 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$1997 \$6905 \$7232 x0_c0_f vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$1998 x0_c0_f_not \$6932 \$6905 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$1999 \$5259 \$6061 \$5995 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2000 \$5996 \$6061 \$5260 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2001 \$5950 \$6061 \$5073 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2002 \$6933 \$6997 \$6063 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2003 \$7451 \$6998 \$6933 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2004 \$6062 \$6905 \$7451 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2005 \$7452 \$6905 \$6063 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2006 \$6934 \$6998 \$7452 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2007 \$5072 \$6061 \$5951 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2008 \$6062 \$6997 \$6934 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2009 x0_c0_b \$6933 \$6905 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$2010 \$6999 \$6934 x0_c0_b vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$2011 x0_c0_b_not \$6933 \$6999 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$2012 \$6905 \$6934 x0_c0_b_not vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$2013 p1 x0_c0_b_not \$6998 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$2014 \$6997 x0_c0_b p1 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$2015 p1_not x0_c0_b_not \$6997 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$2016 \$6998 x0_c0_b p1_not vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$2017 \$5998 a1|b0_p1|b1_p1|b2_p1|b3_p1|b4_p1|b5_p1|b6_p1|b7_p1 b2_c1_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2018 b2_c1 a1|b0_p1|b1_p1|b2_p1|b3_p1|b4_p1|b5_p1|b6_p1|b7_p1 \$5999 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2019 \$7004 \$7238 \$6065 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$2020 \$6064 \$6936 \$7004 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$2021 \$7005 \$7238 \$6064 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$2022 \$6065 \$6936 \$7005 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$2023 \$7006 \$7238 \$7239 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$2024 \$7080 \$6936 \$7006 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$2025 \$6907 \$7238 \$7080 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$2026 \$7239 \$6936 \$6907 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$2027 \$5270 \$6068 \$5998 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2028 \$5999 \$6068 \$5271 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2029 b2_r1_b_not \$6068 \$5077 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$2030 b2_r0_b_not \$7004 \$6070 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$2031 \$7457 \$7005 b2_r0_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$2032 \$6069 \$6907 \$7457 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2033 \$7458 \$6907 \$6070 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2034 b2_r0_b \$7005 \$7458 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2035 \$5076 \$6068 b2_r1_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2036 \$6069 \$7004 b2_r0_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2037 \$7007 b2_r0_b_not \$6907 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$2038 \$7006 b2_r0_b \$7007 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$2039 \$7008 b2_r0_b_not \$7006 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$2040 \$6907 b2_r0_b \$7008 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$2041 p2 \$7008 \$7005 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$2042 \$7004 \$7007 p2 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$2043 p2_not \$7008 \$7004 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$2044 \$7005 \$7007 p2_not vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$2045 \$5956 a1|b0_p1|b1_p1|b2_p1|b3_p1|b4_p1|b5_p1|b6_p1|b7_p1 b2_c1_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2046 b3_c1 a1|b0_p1|b1_p1|b2_p1|b3_p1|b4_p1|b5_p1|b6_p1|b7_p1 \$6000 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2047 \$7011 \$6940 \$6072 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$2048 \$6071 \$6941 \$7011 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$2049 \$7012 \$6940 \$6071 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$2050 \$6072 \$6941 \$7012 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$2051 \$7013 \$6940 \$7242 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$2052 \$7088 \$6941 \$7013 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$2053 \$6908 \$6940 \$7088 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$2054 \$7242 \$6941 \$6908 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$2055 \$5278 \$6075 \$5956 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2056 \$6180 \$7011 \$6940 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2057 \$7461 \$7012 \$6180 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2058 \$6941 \$6908 \$7461 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2059 \$7462 \$6908 \$6940 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2060 \$6416 \$7012 \$7462 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2061 \$6000 \$6075 \$5279 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2062 \$6941 \$7011 \$6416 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2063 b3_r1_b_not \$6075 \$5084 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$2064 b3_r0_b_not \$7011 \$6077 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$2065 \$7463 \$7012 b3_r0_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$2066 \$6076 \$6908 \$7463 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2067 \$7464 \$6908 \$6077 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2068 b3_r0_b \$7012 \$7464 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2069 \$5083 \$6075 b3_r1_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2070 \$6076 \$7011 b3_r0_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2071 \$7014 b3_r0_b_not \$6908 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$2072 \$7013 b3_r0_b \$7014 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$2073 \$7015 b3_r0_b_not \$7013 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$2074 \$6908 b3_r0_b \$7015 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$2075 p3 \$7015 \$7012 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$2076 \$7011 \$7014 p3 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$2077 p3_not \$7015 \$7011 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$2078 \$7012 \$7014 p3_not vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$2079 \$6002 b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b4|b4_q7 b2_c1_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2080 \$6002 a1|b0_p1|b1_p1|b2_p1|b3_p1|b4_p1|b5_p1|b6_p1|b7_p1 b2_c1_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2081 \$6505
+ b2_q0_not|b2_q1_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b4_not|b4_q7_not
+ \$6002 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2082 b4_c1
+ a1_not|b0_p1_not|b1_p1_not|b2_p1_not|b3_p1_not|b4_p1_not|b5_p1_not|b6_p1_not|b7_p1_not
+ \$6505 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2083 \$6506
+ a1_not|b0_p1_not|b1_p1_not|b2_p1_not|b3_p1_not|b4_p1_not|b5_p1_not|b6_p1_not|b7_p1_not
+ b2_c1_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2084 \$6003
+ b2_q0_not|b2_q1_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b4_not|b4_q7_not
+ \$6506 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2085 b4_c1 a1|b0_p1|b1_p1|b2_p1|b3_p1|b4_p1|b5_p1|b6_p1|b7_p1 \$6003 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2086 b4_c1 b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b4|b4_q7 \$6003 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2087 \$7018 \$7248 \$6079 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$2088 \$6078 \$6945 \$7018 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$2089 \$7019 \$7248 \$6078 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$2090 \$6079 \$6945 \$7019 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$2091 \$7020 \$7248 \$7249 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$2092 \$7093 \$6945 \$7020 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$2093 \$6909 \$7248 \$7093 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$2094 \$7249 \$6945 \$6909 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$2095 \$5289 \$6082 \$6002 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2096 \$6188 \$7018 \$7248 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2097 \$7467 \$7019 \$6188 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2098 \$6945 \$6909 \$7467 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2099 \$7468 \$6909 \$7248 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2100 \$6419 \$7019 \$7468 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2101 \$6003 \$6082 \$5290 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2102 \$6945 \$7018 \$6419 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2103 b4_r1_b_not \$6082 \$5089 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$2104 b4_r0_b_not \$7018 \$6084 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$2105 \$7469 \$7019 b4_r0_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$2106 \$6083 \$6909 \$7469 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2107 \$7470 \$6909 \$6084 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2108 b4_r0_b \$7019 \$7470 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2109 \$5088 \$6082 b4_r1_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2110 \$6083 \$7018 b4_r0_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2111 \$7021 b4_r0_b_not \$6909 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$2112 \$7020 b4_r0_b \$7021 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$2113 \$7022 b4_r0_b_not \$7020 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$2114 \$6909 b4_r0_b \$7022 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$2115 p4 \$7022 \$7019 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$2116 \$7018 \$7021 p4 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$2117 p4_not \$7022 \$7018 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$2118 \$7019 \$7021 p4_not vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$2119 \$6005 a1|b0_p1|b1_p1|b2_p1|b3_p1|b4_p1|b5_p1|b6_p1|b7_p1 \$6004 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2120 \$6005 b5|b5_q0|b5_q1|b5_q2|b5_q3|b5_q4|b5_q5|b5_q6|b5_q7 \$6004 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2121 \$6510
+ b5_not|b5_q0_not|b5_q1_not|b5_q2_not|b5_q3_not|b5_q4_not|b5_q5_not|b5_q6_not|b5_q7_not
+ \$6005 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2122 b5_c1
+ a1_not|b0_p1_not|b1_p1_not|b2_p1_not|b3_p1_not|b4_p1_not|b5_p1_not|b6_p1_not|b7_p1_not
+ \$6510 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2123 \$6511
+ a1_not|b0_p1_not|b1_p1_not|b2_p1_not|b3_p1_not|b4_p1_not|b5_p1_not|b6_p1_not|b7_p1_not
+ \$6004 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2124 \$6006
+ b5_not|b5_q0_not|b5_q1_not|b5_q2_not|b5_q3_not|b5_q4_not|b5_q5_not|b5_q6_not|b5_q7_not
+ \$6511 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2125 b5_c1 b5|b5_q0|b5_q1|b5_q2|b5_q3|b5_q4|b5_q5|b5_q6|b5_q7 \$6006 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2126 b5_c1 a1|b0_p1|b1_p1|b2_p1|b3_p1|b4_p1|b5_p1|b6_p1|b7_p1 \$6006 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2127 \$7025 \$7254 \$6086 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$2128 \$6085 \$6949 \$7025 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$2129 \$7026 \$7254 \$6085 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$2130 \$6086 \$6949 \$7026 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$2131 \$7027 \$7254 \$7255 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$2132 \$7098 \$6949 \$7027 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$2133 \$6910 \$7254 \$7098 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$2134 \$7255 \$6949 \$6910 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$2135 \$5299 \$6089 \$6005 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2136 \$6196 \$7025 \$7254 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2137 \$7473 \$7026 \$6196 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2138 \$6949 \$6910 \$7473 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2139 \$7474 \$6910 \$7254 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2140 \$6422 \$7026 \$7474 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2141 \$6006 \$6089 \$5300 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2142 \$6949 \$7025 \$6422 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2143 b5_r1_b_not \$6089 \$5094 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$2144 b5_r0_b_not \$7025 \$6091 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$2145 \$7475 \$7026 b5_r0_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$2146 \$6090 \$6910 \$7475 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2147 \$7476 \$6910 \$6091 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2148 b5_r0_b \$7026 \$7476 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2149 \$5093 \$6089 b5_r1_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2150 \$6090 \$7025 b5_r0_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2151 \$7028 b5_r0_b_not \$6910 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$2152 \$7027 b5_r0_b \$7028 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$2153 \$7029 b5_r0_b_not \$7027 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$2154 \$6910 b5_r0_b \$7029 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$2155 p5 \$7029 \$7026 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$2156 \$7025 \$7028 p5 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$2157 p5_not \$7029 \$7025 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$2158 \$7026 \$7028 p5_not vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$2159 \$6008 a1|b0_p1|b1_p1|b2_p1|b3_p1|b4_p1|b5_p1|b6_p1|b7_p1 b6_c1_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2160 b6_c1 a1|b0_p1|b1_p1|b2_p1|b3_p1|b4_p1|b5_p1|b6_p1|b7_p1 \$6009 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2161 \$7032 \$7261 \$6093 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$2162 \$6092 \$6954 \$7032 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$2163 \$7033 \$7261 \$6092 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$2164 \$6093 \$6954 \$7033 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$2165 \$7034 \$7261 \$7262 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$2166 \$7103 \$6954 \$7034 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$2167 \$6911 \$7261 \$7103 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$2168 \$7262 \$6954 \$6911 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$2169 \$5308 \$6096 \$6008 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2170 \$6203 \$7032 \$7261 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2171 \$7479 \$7033 \$6203 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2172 \$6954 \$6911 \$7479 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2173 \$7480 \$6911 \$7261 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2174 \$6425 \$7033 \$7480 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2175 \$6009 \$6096 \$5309 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2176 \$6954 \$7032 \$6425 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2177 b6_r1_b_not \$6096 \$5099 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$2178 b6_r0_b_not \$7032 \$6098 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$2179 \$7481 \$7033 b6_r0_b_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$2180 \$6097 \$6911 \$7481 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2181 \$7482 \$6911 \$6098 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2182 b6_r0_b \$7033 \$7482 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2183 \$5098 \$6096 b6_r1_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2184 \$6097 \$7032 b6_r0_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2185 \$7035 b6_r0_b_not \$6911 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$2186 \$7034 b6_r0_b \$7035 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$2187 \$7036 b6_r0_b_not \$7034 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$2188 \$6911 b6_r0_b \$7036 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$2189 p6 \$7036 \$7033 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$2190 \$7032 \$7035 p6 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$2191 p6_not \$7036 \$7032 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$2192 \$7033 \$7035 p6_not vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$2193 \$6011 a1|b0_p1|b1_p1|b2_p1|b3_p1|b4_p1|b5_p1|b6_p1|b7_p1 \$6010 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2194 b6_c1 a1|b0_p1|b1_p1|b2_p1|b3_p1|b4_p1|b5_p1|b6_p1|b7_p1 \$6012 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2195 \$7039 \$7267 \$6100 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$2196 \$6099 \$6958 \$7039 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$2197 \$7040 \$7267 \$6099 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$2198 \$6100 \$6958 \$7040 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$2199 \$7041 \$7267 \$7268 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$2200 \$7108 \$6958 \$7041 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$2201 \$6912 \$7267 \$7108 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$2202 \$7268 \$6958 \$6912 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$2203 \$5318 \$6103 \$6011 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2204 \$6211 \$7039 \$7267 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2205 \$7485 \$7040 \$6211 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2206 \$6958 \$6912 \$7485 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2207 \$7486 \$6912 \$7267 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2208 \$6427 \$7040 \$7486 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2209 \$6012 \$6103 \$5319 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2210 \$6958 \$7039 \$6427 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2211 \$5970 \$6103 \$5104 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2212 \$6960 \$7039 \$6105 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2213 \$7487 \$7040 \$6960 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2214 \$6104 \$6912 \$7487 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2215 \$7488 \$6912 \$6105 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2216 \$6961 \$7040 \$7488 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2217 \$5103 \$6103 \$5971 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2218 \$6104 \$7039 \$6961 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2219 \$7042 \$6960 \$6912 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P
+ AD=0.6669P PS=3.45U PD=3.55U
M$2220 \$7041 \$6961 \$7042 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P
+ AD=0.60515P PS=3.55U PD=3.45U
M$2221 \$7043 \$6960 \$7041 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$2222 \$6912 \$6961 \$7043 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$2223 p7 \$7043 \$7040 vdd pfet_03v3 L=0.5U W=1.235U AS=0.60515P AD=0.6669P
+ PS=3.45U PD=3.55U
M$2224 \$7039 \$7042 p7 vdd pfet_03v3 L=0.5U W=1.235U AS=0.6669P AD=0.60515P
+ PS=3.55U PD=3.45U
M$2225 p7_not \$7043 \$7039 vdd pfet_03v3 L=0.5U W=1.235U AS=0.648375P
+ AD=0.60515P PS=3.52U PD=3.45U
M$2226 \$7040 \$7042 p7_not vdd pfet_03v3 L=0.5U W=1.235U AS=0.6422P
+ AD=0.70395P PS=3.51U PD=3.61U
M$2227 \$6929 a0|b0_p0|b1_p0|b2_p0|b3_p0|b4_p0|b5_p0|b6_p0|b7_p0 b1_c0_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2228 b1_c0 a0|b0_p0|b1_p0|b2_p0|b3_p0|b4_p0|b5_p0|b6_p0|b7_p0 \$6930 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2229 p0_not b0|b0_q0|b0_q1|b0_q2|b0_q3|b0_q4|b0_q5|b0_q6|b0_q7 b0_c0_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2230 p0_not a0|b0_p0|b1_p0|b2_p0|b3_p0|b4_p0|b5_p0|b6_p0|b7_p0 b0_c0_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2231 \$7232 b0|b0_q0|b0_q1|b0_q2|b0_q3|b0_q4|b0_q5|b0_q6|b0_q7 b0_c1_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2232 \$7232 a1|b0_p1|b1_p1|b2_p1|b3_p1|b4_p1|b5_p1|b6_p1|b7_p1 b0_c1_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2233 \$7884
+ b0_not|b0_q0_not|b0_q1_not|b0_q3_not|b0_q4_not|b0_q5_not|b0_q6_not|b0_q7_not|b1_q2_not
+ p0_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2234 \$7447
+ b0_not|b0_q0_not|b0_q1_not|b0_q3_not|b0_q4_not|b0_q5_not|b0_q6_not|b0_q7_not|b1_q2_not
+ \$7232 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2235 b0_c0
+ a0_not|b0_p0_not|b1_p0_not|b2_p0_not|b3_p0_not|b5_p0_not|b6_p0_not|b7_p0_not
+ \$7884 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2236 b0_c1
+ a1_not|b0_p1_not|b1_p1_not|b2_p1_not|b3_p1_not|b4_p1_not|b5_p1_not|b6_p1_not|b7_p1_not
+ \$7447 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2237 \$7885
+ a0_not|b0_p0_not|b1_p0_not|b2_p0_not|b3_p0_not|b5_p0_not|b6_p0_not|b7_p0_not
+ b0_c0_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2238 \$7448
+ a1_not|b0_p1_not|b1_p1_not|b2_p1_not|b3_p1_not|b4_p1_not|b5_p1_not|b6_p1_not|b7_p1_not
+ b0_c1_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2239 p0
+ b0_not|b0_q0_not|b0_q1_not|b0_q3_not|b0_q4_not|b0_q5_not|b0_q6_not|b0_q7_not|b1_q2_not
+ \$7885 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2240 \$6932
+ b0_not|b0_q0_not|b0_q1_not|b0_q3_not|b0_q4_not|b0_q5_not|b0_q6_not|b0_q7_not|b1_q2_not
+ \$7448 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2241 b0_c0 a0|b0_p0|b1_p0|b2_p0|b3_p0|b4_p0|b5_p0|b6_p0|b7_p0 p0 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2242 b0_c0 b0|b0_q0|b0_q1|b0_q2|b0_q3|b0_q4|b0_q5|b0_q6|b0_q7 p0 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2243 b0_c1 b0|b0_q0|b0_q1|b0_q2|b0_q3|b0_q4|b0_q5|b0_q6|b0_q7 \$6932 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2244 b0_c1 a1|b0_p1|b1_p1|b2_p1|b3_p1|b4_p1|b5_p1|b6_p1|b7_p1 \$6932 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2245 \$6164 \$6999 \$7232 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2246 \$6164 \$6997 \$7232 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2247 \$7449 \$6998 \$6164 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2248 \$6932 \$6905 \$7449 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2249 \$7450 \$6905 \$7232 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2250 \$6411 \$6998 \$7450 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2251 \$6932 \$6997 \$6411 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2252 \$6932 \$6999 \$6411 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2253 \$6933 \$6999 \$6063 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2254 \$6062 \$6999 \$6934 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2255 \$7238 b2|b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7 b2_c0_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2256 \$7238 a0|b0_p0|b1_p0|b2_p0|b3_p0|b4_p0|b5_p0|b6_p0|b7_p0 b2_c0_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2257 \$7453
+ b2_not|b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not
+ \$7238 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2258 b2_c0
+ a0_not|b0_p0_not|b1_p0_not|b2_p0_not|b3_p0_not|b5_p0_not|b6_p0_not|b7_p0_not
+ \$7453 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2259 \$7454
+ a0_not|b0_p0_not|b1_p0_not|b2_p0_not|b3_p0_not|b5_p0_not|b6_p0_not|b7_p0_not
+ b2_c0_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2260 \$6936
+ b2_not|b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not
+ \$7454 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2261 b2_c0 b2|b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7 \$6936 vdd pfet_03v3
+ L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2262 b2_c0 a0|b0_p0|b1_p0|b2_p0|b3_p0|b4_p0|b5_p0|b6_p0|b7_p0 \$6936 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2263 \$6172 \$7006 \$7238 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2264 \$6172 \$7004 \$7238 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2265 \$7455 \$7005 \$6172 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2266 \$6936 \$6907 \$7455 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2267 \$7456 \$6907 \$7238 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2268 \$6413 \$7005 \$7456 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2269 \$6936 \$7004 \$6413 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2270 \$6936 \$7006 \$6413 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2271 b2_r0_b_not \$7006 \$6070 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$2272 \$6069 \$7006 b2_r0_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2273 \$6940 a0|b0_p0|b1_p0|b2_p0|b3_p0|b4_p0|b5_p0|b6_p0|b7_p0 b2_c0_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2274 \$6940
+ b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b3|b3_q0|b3_q1|b3_q2|b3_q3|b3_q4|b3_q5|b3_q6|b3_q7
+ b2_c0_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2275 \$7459
+ b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b3_not|b3_q0_not|b3_q1_not|b3_q2_not|b3_q3_not|b3_q4_not|b3_q5_not|b3_q6_not|b3_q7_not
+ \$6940 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2276 b2_c0
+ a0_not|b0_p0_not|b1_p0_not|b2_p0_not|b3_p0_not|b5_p0_not|b6_p0_not|b7_p0_not
+ \$7459 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2277 \$7460
+ a0_not|b0_p0_not|b1_p0_not|b2_p0_not|b3_p0_not|b5_p0_not|b6_p0_not|b7_p0_not
+ b2_c0_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2278 \$6941
+ b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b3_not|b3_q0_not|b3_q1_not|b3_q2_not|b3_q3_not|b3_q4_not|b3_q5_not|b3_q6_not|b3_q7_not
+ \$7460 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2279 b2_c0 a0|b0_p0|b1_p0|b2_p0|b3_p0|b4_p0|b5_p0|b6_p0|b7_p0 \$6941 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2280 b2_c0
+ b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b3|b3_q0|b3_q1|b3_q2|b3_q3|b3_q4|b3_q5|b3_q6|b3_q7
+ \$6941 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2281 \$6180 \$7013 \$6940 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2282 \$6941 \$7013 \$6416 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2283 b3_r0_b_not \$7013 \$6077 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$2284 \$6076 \$7013 b3_r0_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2285 \$7248 a0|b0_p0|b1_p0|b2_p0|b3_p0|b4_p0|b5_p0|b6_p0|b7_p0 b2_c0_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2286 \$7248 b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b4|b4_q7 b2_c0_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2287 \$7465
+ b2_q0_not|b2_q1_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b4_not|b4_q7_not
+ \$7248 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2288 b2_c0
+ a0_not|b0_p0_not|b1_p0_not|b2_p0_not|b3_p0_not|b5_p0_not|b6_p0_not|b7_p0_not
+ \$7465 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2289 \$7466
+ a0_not|b0_p0_not|b1_p0_not|b2_p0_not|b3_p0_not|b5_p0_not|b6_p0_not|b7_p0_not
+ b2_c0_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2290 \$6945
+ b2_q0_not|b2_q1_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b4_not|b4_q7_not
+ \$7466 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2291 b2_c0 a0|b0_p0|b1_p0|b2_p0|b3_p0|b4_p0|b5_p0|b6_p0|b7_p0 \$6945 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2292 b2_c0 b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b4|b4_q7 \$6945 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2293 \$6188 \$7020 \$7248 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2294 \$6945 \$7020 \$6419 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2295 b4_r0_b_not \$7020 \$6084 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$2296 \$6083 \$7020 b4_r0_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2297 \$7254 a0|b0_p0|b1_p0|b2_p0|b3_p0|b4_p0|b5_p0|b6_p0|b7_p0 \$6948 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2298 \$7254 b5|b5_q0|b5_q1|b5_q2|b5_q3|b5_q4|b5_q5|b5_q6|b5_q7 \$6948 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2299 \$7471
+ b5_not|b5_q0_not|b5_q1_not|b5_q2_not|b5_q3_not|b5_q4_not|b5_q5_not|b5_q6_not|b5_q7_not
+ \$7254 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2300 \$6950
+ a0_not|b0_p0_not|b1_p0_not|b2_p0_not|b3_p0_not|b5_p0_not|b6_p0_not|b7_p0_not
+ \$7471 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2301 \$7472
+ a0_not|b0_p0_not|b1_p0_not|b2_p0_not|b3_p0_not|b5_p0_not|b6_p0_not|b7_p0_not
+ \$6948 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2302 \$6949
+ b5_not|b5_q0_not|b5_q1_not|b5_q2_not|b5_q3_not|b5_q4_not|b5_q5_not|b5_q6_not|b5_q7_not
+ \$7472 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2303 \$6950 a0|b0_p0|b1_p0|b2_p0|b3_p0|b4_p0|b5_p0|b6_p0|b7_p0 \$6949 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2304 \$6950 b5|b5_q0|b5_q1|b5_q2|b5_q3|b5_q4|b5_q5|b5_q6|b5_q7 \$6949 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2305 \$6196 \$7027 \$7254 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2306 \$6949 \$7027 \$6422 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2307 b5_r0_b_not \$7027 \$6091 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$2308 \$6090 \$7027 b5_r0_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2309 \$7261 b6|b6_q0|b6_q1|b6_q2|b6_q3|b6_q4|b6_q5|b6_q6|b6_q7 b6_c0_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2310 \$7261 a0|b0_p0|b1_p0|b2_p0|b3_p0|b4_p0|b5_p0|b6_p0|b7_p0 b6_c0_not vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2311 \$7477
+ b6_not|b6_q0_not|b6_q1_not|b6_q2_not|b6_q3_not|b6_q4_not|b6_q5_not|b6_q6_not|b6_q7_not
+ \$7261 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2312 b6_c0
+ a0_not|b0_p0_not|b1_p0_not|b2_p0_not|b3_p0_not|b5_p0_not|b6_p0_not|b7_p0_not
+ \$7477 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2313 \$7478
+ a0_not|b0_p0_not|b1_p0_not|b2_p0_not|b3_p0_not|b5_p0_not|b6_p0_not|b7_p0_not
+ b6_c0_not vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2314 \$6954
+ b6_not|b6_q0_not|b6_q1_not|b6_q2_not|b6_q3_not|b6_q4_not|b6_q5_not|b6_q6_not|b6_q7_not
+ \$7478 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2315 b6_c0 a0|b0_p0|b1_p0|b2_p0|b3_p0|b4_p0|b5_p0|b6_p0|b7_p0 \$6954 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2316 b6_c0 b6|b6_q0|b6_q1|b6_q2|b6_q3|b6_q4|b6_q5|b6_q6|b6_q7 \$6954 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2317 \$6203 \$7034 \$7261 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2318 \$6954 \$7034 \$6425 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2319 b6_r0_b_not \$7034 \$6098 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P
+ AD=0.273P PS=2.14U PD=2.14U
M$2320 \$6097 \$7034 b6_r0_b vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2321 \$7267 b1_q3|b7|b7_q0|b7_q1|b7_q2|b7_q4|b7_q5|b7_q6|b7_q7 \$6957 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2322 \$7267 a0|b0_p0|b1_p0|b2_p0|b3_p0|b4_p0|b5_p0|b6_p0|b7_p0 \$6957 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2323 \$7483
+ b7_not|b7_q0_not|b7_q1_not|b7_q2_not|b7_q3_not|b7_q4_not|b7_q5_not|b7_q6_not|b7_q7_not
+ \$7267 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2324 \$6959
+ a0_not|b0_p0_not|b1_p0_not|b2_p0_not|b3_p0_not|b5_p0_not|b6_p0_not|b7_p0_not
+ \$7483 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2325 \$7484
+ a0_not|b0_p0_not|b1_p0_not|b2_p0_not|b3_p0_not|b5_p0_not|b6_p0_not|b7_p0_not
+ \$6957 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2326 \$6958
+ b7_not|b7_q0_not|b7_q1_not|b7_q2_not|b7_q3_not|b7_q4_not|b7_q5_not|b7_q6_not|b7_q7_not
+ \$7484 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2327 \$6959 a0|b0_p0|b1_p0|b2_p0|b3_p0|b4_p0|b5_p0|b6_p0|b7_p0 \$6958 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2328 \$6959 b1_q3|b7|b7_q0|b7_q1|b7_q2|b7_q4|b7_q5|b7_q6|b7_q7 \$6958 vdd
+ pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P PS=2.14U PD=2.14U
M$2329 \$6211 \$7041 \$7267 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2330 \$6958 \$7041 \$6427 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2331 \$6960 \$7041 \$6105 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2332 \$6104 \$7041 \$6961 vdd pfet_03v3 L=0.28U W=0.42U AS=0.273P AD=0.273P
+ PS=2.14U PD=2.14U
M$2333 x2_b0_f \$80 \$15 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2334 x2_b0_f_not \$80 \$17 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2335 \$15 \$166 x2_b0_f_not vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$2336 \$17 \$166 x2_b0_f vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2337 x3_b0_f \$82 \$34 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2338 x4_b0_f \$84 \$36 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2339 x5_b0_f \$86 \$38 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2340 x6_b0_f \$88 p15 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2341 x0_b0_f \$76 \$27 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2342 x0_b0_f_not \$76 \$28 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2343 x1_b0_f \$78 \$30 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2344 x1_b0_f_not \$78 \$31 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2345 x3_b0_f_not \$82 \$19 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2346 x4_b0_f_not \$84 \$21 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2347 x5_b0_f_not \$86 \$23 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2348 x6_b0_f_not \$88 p15_not vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2349 \$220
+ a7_not|b0_p7_not|b1_p7_not|b2_p7_not|b4_p7_not|b5_p7_not|b6_p7_not|b7_p7_not
+ b1_c7_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2350 b1_c7
+ a7_not|b0_p7_not|b1_p7_not|b2_p7_not|b4_p7_not|b5_p7_not|b6_p7_not|b7_p7_not
+ \$151 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2351 \$27 \$152 x0_b0_f_not vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$2352 \$28 \$152 x0_b0_f vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2353 \$30 \$159 x1_b0_f_not vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$2354 \$31 \$159 x1_b0_f vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2355 b3_r7_b_not \$145 \$80 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2356 \$166 \$145 b3_r7_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2357 \$34 \$173 x3_b0_f_not vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$2358 \$19 \$173 x3_b0_f vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2359 \$36 \$180 x4_b0_f_not vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$2360 \$21 \$180 x4_b0_f vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2361 \$38 \$187 x5_b0_f_not vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$2362 \$23 \$187 x5_b0_f vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2363 p15 \$194 x6_b0_f_not vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$2364 p15_not \$194 x6_b0_f vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2365 \$80 \$145 \$163 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2366 \$165 \$145 \$166 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2367 b4_r7_b_not \$146 \$82 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2368 \$173 \$146 b4_r7_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2369 b5_r7_b_not \$147 \$84 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2370 \$180 \$147 b5_r7_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2371 b6_r7_b_not \$148 \$86 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2372 \$187 \$148 b6_r7_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2373 \$195 \$149 \$88 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2374 \$194 \$149 \$196 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2375 \$76 \$142 x0_a7_f_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2376 x0_a7_f \$142 \$152 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2377 x0_a7_b_not \$142 \$76 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2378 \$152 \$142 x0_a7_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2379 \$78 \$143 \$156 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2380 \$158 \$143 \$159 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2381 b2_r7_b_not \$143 \$78 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2382 \$159 \$143 b2_r7_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2383 \$82 \$146 \$170 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2384 \$172 \$146 \$173 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2385 \$84 \$147 \$177 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2386 \$179 \$147 \$180 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2387 \$86 \$148 \$184 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2388 \$186 \$148 \$187 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2389 \$88 \$149 \$191 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2390 \$193 \$149 \$194 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2391 \$156
+ a7_not|b0_p7_not|b1_p7_not|b2_p7_not|b4_p7_not|b5_p7_not|b6_p7_not|b7_p7_not
+ b2_c7_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2392 b2_c7
+ a7_not|b0_p7_not|b1_p7_not|b2_p7_not|b4_p7_not|b5_p7_not|b6_p7_not|b7_p7_not
+ \$158 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2393 \$163 b2_p7_not|b3_p7_not b3_c7_not vss nfet_03v3 L=0.28U W=0.42U
+ AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2394 b3_c7 b2_p7_not|b3_p7_not \$165 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2395 \$287 \$165 \$30 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2396 \$31 \$163 \$287 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2397 \$30 \$163 \$289 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P AD=0.6925P
+ PS=3.74U PD=3.77U
M$2398 \$288 \$165 \$223 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2399 \$451 \$163 \$288 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2400 \$223 \$163 \$145 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P AD=0.6925P
+ PS=3.74U PD=3.77U
M$2401 \$290 b3_r7_b \$145 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2402 \$288 b3_r7_b_not \$290 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2403 \$291 b3_r7_b \$288 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2404 \$145 b3_r7_b_not \$291 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2405 \$292 \$290 \$289 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2406 \$287 \$291 \$292 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2407 \$293 \$290 \$287 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2408 \$289 \$291 \$293 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P AD=0.6925P
+ PS=3.74U PD=3.77U
M$2409 \$170
+ a7_not|b0_p7_not|b1_p7_not|b2_p7_not|b4_p7_not|b5_p7_not|b6_p7_not|b7_p7_not
+ b4_c7_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2410 b4_c7
+ a7_not|b0_p7_not|b1_p7_not|b2_p7_not|b4_p7_not|b5_p7_not|b6_p7_not|b7_p7_not
+ \$172 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2411 \$297 b4_r7_b_not \$298 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2412 \$295 \$299 \$300 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2413 \$177
+ a7_not|b0_p7_not|b1_p7_not|b2_p7_not|b4_p7_not|b5_p7_not|b6_p7_not|b7_p7_not
+ b5_c7_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2414 b5_c7
+ a7_not|b0_p7_not|b1_p7_not|b2_p7_not|b4_p7_not|b5_p7_not|b6_p7_not|b7_p7_not
+ \$179 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2415 \$305 b5_r7_b_not \$306 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2416 \$303 \$307 \$308 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2417 \$184
+ a7_not|b0_p7_not|b1_p7_not|b2_p7_not|b4_p7_not|b5_p7_not|b6_p7_not|b7_p7_not
+ b6_c7_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2418 b6_c7
+ a7_not|b0_p7_not|b1_p7_not|b2_p7_not|b4_p7_not|b5_p7_not|b6_p7_not|b7_p7_not
+ \$186 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2419 \$313 b6_r7_b_not \$314 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2420 \$311 \$315 \$316 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2421 \$191
+ a7_not|b0_p7_not|b1_p7_not|b2_p7_not|b4_p7_not|b5_p7_not|b6_p7_not|b7_p7_not
+ b6_c7_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2422 b6_c7
+ a7_not|b0_p7_not|b1_p7_not|b2_p7_not|b4_p7_not|b5_p7_not|b6_p7_not|b7_p7_not
+ \$193 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2423 \$321 \$195 \$322 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2424 \$319 \$323 p14 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P AD=0.657975P
+ PS=3.88U PD=3.76U
M$2425 \$151 x0_a7_f_not \$271 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2426 \$220 x0_a7_f_not \$272 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2427 \$608 x0_a7_f_not \$273 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2428 \$221 x0_a7_f_not \$142 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2429 \$273 x0_a7_b_not \$274 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2430 \$142 x0_a7_b_not \$275 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2431 \$271 \$275 \$276 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2432 \$272 \$275 \$277 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P AD=0.6925P
+ PS=3.74U PD=3.77U
M$2433 \$28 \$156 \$279 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2434 \$27 \$156 \$280 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P AD=0.6925P
+ PS=3.74U PD=3.77U
M$2435 \$613 \$156 \$281 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2436 \$222 \$156 \$143 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P AD=0.6925P
+ PS=3.74U PD=3.77U
M$2437 \$281 b2_r7_b_not \$282 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2438 \$143 b2_r7_b_not \$283 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2439 \$279 \$283 \$284 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2440 \$280 \$283 \$285 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P AD=0.6925P
+ PS=3.74U PD=3.77U
M$2441 \$289 \$165 \$31 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P AD=0.64155P
+ PS=3.68U PD=3.67U
M$2442 \$145 \$165 \$451 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2443 \$295 \$172 \$15 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2444 \$17 \$170 \$295 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2445 \$15 \$170 \$296 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P AD=0.6925P
+ PS=3.74U PD=3.77U
M$2446 \$297 \$172 \$224 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2447 \$622 \$170 \$297 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2448 \$224 \$170 \$146 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P AD=0.6925P
+ PS=3.74U PD=3.77U
M$2449 \$298 b4_r7_b \$146 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2450 \$299 b4_r7_b \$297 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2451 \$146 b4_r7_b_not \$299 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2452 \$300 \$298 \$296 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2453 \$301 \$298 \$295 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2454 \$296 \$299 \$301 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P AD=0.6925P
+ PS=3.74U PD=3.77U
M$2455 \$303 \$179 \$34 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2456 \$19 \$177 \$303 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2457 \$34 \$177 \$304 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P AD=0.6925P
+ PS=3.74U PD=3.77U
M$2458 \$305 \$179 \$225 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2459 \$627 \$177 \$305 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2460 \$225 \$177 \$147 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P AD=0.6925P
+ PS=3.74U PD=3.77U
M$2461 \$306 b5_r7_b \$147 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2462 \$307 b5_r7_b \$305 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2463 \$147 b5_r7_b_not \$307 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2464 \$308 \$306 \$304 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2465 \$309 \$306 \$303 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2466 \$304 \$307 \$309 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P AD=0.6925P
+ PS=3.74U PD=3.77U
M$2467 \$311 \$186 \$36 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2468 \$21 \$184 \$311 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2469 \$36 \$184 \$312 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P AD=0.6925P
+ PS=3.74U PD=3.77U
M$2470 \$313 \$186 \$226 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2471 \$632 \$184 \$313 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2472 \$226 \$184 \$148 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P AD=0.6925P
+ PS=3.74U PD=3.77U
M$2473 \$314 b6_r7_b \$148 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2474 \$315 b6_r7_b \$313 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2475 \$148 b6_r7_b_not \$315 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2476 \$316 \$314 \$312 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2477 \$317 \$314 \$311 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2478 \$312 \$315 \$317 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P AD=0.6925P
+ PS=3.74U PD=3.77U
M$2479 \$319 \$193 \$38 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2480 \$23 \$191 \$319 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2481 \$38 \$191 \$320 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P AD=0.6925P
+ PS=3.74U PD=3.77U
M$2482 \$321 \$193 \$227 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2483 \$637 \$191 \$321 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2484 \$227 \$191 \$149 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P AD=0.6925P
+ PS=3.74U PD=3.77U
M$2485 \$322 \$196 \$149 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2486 \$323 \$196 \$321 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2487 \$149 \$195 \$323 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P AD=0.6925P
+ PS=3.74U PD=3.77U
M$2488 p14 \$322 \$320 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2489 p14_not \$322 \$319 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2490 \$320 \$323 p14_not vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2491 \$220
+ b1_not|b1_q0_not|b1_q1_not|b1_q2_not|b1_q3_not|b1_q4_not|b1_q5_not|b1_q6_not|b1_q7_not
+ b1_c7_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2492 \$436 a7|b0_p7|b1_p7|b2_p7|b3_p7|b4_p7|b5_p7|b6_p7|b7_p7 \$220 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2493 b1_c7 b1|b1_q0|b1_q1|b1_q2|b1_q3|b1_q4|b1_q5|b1_q6|b1_q7 \$436 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2494 \$438 b1|b1_q0|b1_q1|b1_q2|b1_q3|b1_q4|b1_q5|b1_q6|b1_q7 b1_c7_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2495 \$151 a7|b0_p7|b1_p7|b2_p7|b3_p7|b4_p7|b5_p7|b6_p7|b7_p7 \$438 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2496 b1_c7
+ b1_not|b1_q0_not|b1_q1_not|b1_q2_not|b1_q3_not|b1_q4_not|b1_q5_not|b1_q6_not|b1_q7_not
+ \$151 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2497 \$271 x0_a7_f \$220 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2498 \$272 x0_a7_f \$151 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2499 \$273 x0_a7_f \$221 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2500 \$142 x0_a7_f \$608 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2501 \$76 \$272 x0_a7_f_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2502 \$439 \$273 \$76 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2503 x0_a7_f \$271 \$439 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2504 \$440 \$271 x0_a7_f_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2505 \$152 \$273 \$440 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2506 x0_a7_f \$272 \$152 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2507 x0_a7_b_not \$272 \$76 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2508 \$441 \$273 x0_a7_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2509 \$152 \$271 \$441 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2510 \$442 \$271 \$76 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2511 x0_a7_b \$273 \$442 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2512 \$152 \$272 x0_a7_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2513 \$274 x0_a7_b \$142 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2514 \$275 x0_a7_b \$273 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2515 \$276 \$274 \$272 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2516 \$277 \$274 \$271 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2517 \$279 \$158 \$27 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2518 \$280 \$158 \$28 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P AD=0.64155P
+ PS=3.68U PD=3.67U
M$2519 \$281 \$158 \$222 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2520 \$143 \$158 \$613 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2521 \$78 \$280 \$156 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2522 \$445 \$281 \$78 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2523 \$158 \$279 \$445 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2524 \$446 \$279 \$156 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2525 \$159 \$281 \$446 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2526 \$158 \$280 \$159 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2527 b2_r7_b_not \$280 \$78 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2528 \$447 \$281 b2_r7_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2529 \$159 \$279 \$447 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2530 \$448 \$279 \$78 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2531 b2_r7_b \$281 \$448 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2532 \$159 \$280 b2_r7_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2533 \$282 b2_r7_b \$143 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2534 \$283 b2_r7_b \$281 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2535 \$284 \$282 \$280 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2536 \$285 \$282 \$279 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2537 \$163
+ b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b3_not|b3_q0_not|b3_q1_not|b3_q2_not|b3_q3_not|b3_q4_not|b3_q5_not|b3_q6_not|b3_q7_not
+ b3_c7_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2538 \$449 a7|b0_p7|b1_p7|b2_p7|b3_p7|b4_p7|b5_p7|b6_p7|b7_p7 \$163 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2539 b3_c7
+ b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b3|b3_q0|b3_q1|b3_q2|b3_q3|b3_q4|b3_q5|b3_q6|b3_q7
+ \$449 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2540 \$450
+ b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b3|b3_q0|b3_q1|b3_q2|b3_q3|b3_q4|b3_q5|b3_q6|b3_q7
+ b3_c7_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2541 \$165 a7|b0_p7|b1_p7|b2_p7|b3_p7|b4_p7|b5_p7|b6_p7|b7_p7 \$450 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2542 b3_c7
+ b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b3_not|b3_q0_not|b3_q1_not|b3_q2_not|b3_q3_not|b3_q4_not|b3_q5_not|b3_q6_not|b3_q7_not
+ \$165 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2543 \$80 \$289 \$163 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2544 \$452 \$288 \$80 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2545 \$165 \$287 \$452 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2546 \$453 \$287 \$163 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2547 \$166 \$288 \$453 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2548 \$165 \$289 \$166 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2549 b3_r7_b_not \$289 \$80 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2550 \$454 \$288 b3_r7_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2551 \$166 \$287 \$454 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2552 \$455 \$287 \$80 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2553 b3_r7_b \$288 \$455 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2554 \$166 \$289 b3_r7_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2555 \$296 \$172 \$17 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P AD=0.64155P
+ PS=3.68U PD=3.67U
M$2556 \$146 \$172 \$622 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2557 \$82 \$296 \$170 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2558 \$458 \$297 \$82 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2559 \$172 \$295 \$458 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2560 \$459 \$295 \$170 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2561 \$173 \$297 \$459 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2562 \$172 \$296 \$173 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2563 b4_r7_b_not \$296 \$82 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2564 \$460 \$297 b4_r7_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2565 \$173 \$295 \$460 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2566 \$461 \$295 \$82 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2567 b4_r7_b \$297 \$461 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2568 \$173 \$296 b4_r7_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2569 \$304 \$179 \$19 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P AD=0.64155P
+ PS=3.68U PD=3.67U
M$2570 \$147 \$179 \$627 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2571 \$84 \$304 \$177 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2572 \$464 \$305 \$84 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2573 \$179 \$303 \$464 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2574 \$465 \$303 \$177 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2575 \$180 \$305 \$465 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2576 \$179 \$304 \$180 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2577 b5_r7_b_not \$304 \$84 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2578 \$466 \$305 b5_r7_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2579 \$180 \$303 \$466 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2580 \$467 \$303 \$84 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2581 b5_r7_b \$305 \$467 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2582 \$180 \$304 b5_r7_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2583 \$312 \$186 \$21 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P AD=0.64155P
+ PS=3.68U PD=3.67U
M$2584 \$148 \$186 \$632 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2585 \$86 \$312 \$184 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2586 \$470 \$313 \$86 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2587 \$186 \$311 \$470 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2588 \$471 \$311 \$184 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2589 \$187 \$313 \$471 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2590 \$186 \$312 \$187 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2591 b6_r7_b_not \$312 \$86 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2592 \$472 \$313 b6_r7_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2593 \$187 \$311 \$472 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2594 \$473 \$311 \$86 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2595 b6_r7_b \$313 \$473 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2596 \$187 \$312 b6_r7_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2597 \$320 \$193 \$23 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P AD=0.64155P
+ PS=3.68U PD=3.67U
M$2598 \$149 \$193 \$637 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2599 \$88 \$320 \$191 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2600 \$476 \$321 \$88 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2601 \$193 \$319 \$476 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2602 \$477 \$319 \$191 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2603 \$194 \$321 \$477 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2604 \$193 \$320 \$194 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2605 \$195 \$320 \$88 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2606 \$478 \$321 \$195 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2607 \$194 \$319 \$478 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2608 \$479 \$319 \$88 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2609 \$196 \$321 \$479 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2610 \$194 \$320 \$196 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2611 \$1397
+ a6_not|b0_p6_not|b1_p6_not|b3_p6_not|b4_p6_not|b5_p6_not|b6_p6_not|b7_p6_not
+ b1_c6_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2612 b1_c6
+ a6_not|b0_p6_not|b1_p6_not|b3_p6_not|b4_p6_not|b5_p6_not|b6_p6_not|b7_p6_not
+ \$1107 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2613 \$1110
+ a7_not|b0_p7_not|b1_p7_not|b2_p7_not|b4_p7_not|b5_p7_not|b6_p7_not|b7_p7_not
+ b0_c7_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2614 b0_c7
+ a7_not|b0_p7_not|b1_p7_not|b2_p7_not|b4_p7_not|b5_p7_not|b6_p7_not|b7_p7_not
+ \$1112 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2615 \$221 \$725 \$1110 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2616 \$1112 \$725 \$608 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2617 b0_r7_b_not \$725 \$275 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2618 \$274 \$725 b0_r7_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2619 \$156
+ b2_not|b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not
+ b2_c7_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2620 \$1117
+ a6_not|b0_p6_not|b1_p6_not|b3_p6_not|b4_p6_not|b5_p6_not|b6_p6_not|b7_p6_not
+ b2_c6_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2621 \$443 a7|b0_p7|b1_p7|b2_p7|b3_p7|b4_p7|b5_p7|b6_p7|b7_p7 \$156 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2622 b2_c7 b2|b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7 \$443 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2623 \$444 b2|b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7 b2_c7_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2624 \$158 a7|b0_p7|b1_p7|b2_p7|b3_p7|b4_p7|b5_p7|b6_p7|b7_p7 \$444 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2625 b2_c7
+ b2_not|b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not
+ \$158 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2626 b2_c6
+ a6_not|b0_p6_not|b1_p6_not|b3_p6_not|b4_p6_not|b5_p6_not|b6_p6_not|b7_p6_not
+ \$1119 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2627 \$222 \$727 \$1117 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2628 \$1119 \$727 \$613 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2629 b2_r6_b_not \$727 \$283 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2630 \$282 \$727 b2_r6_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2631 \$1123
+ a6_not|b0_p6_not|b1_p6_not|b3_p6_not|b4_p6_not|b5_p6_not|b6_p6_not|b7_p6_not
+ b3_c6_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2632 b3_c6
+ a6_not|b0_p6_not|b1_p6_not|b3_p6_not|b4_p6_not|b5_p6_not|b6_p6_not|b7_p6_not
+ \$1125 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2633 \$223 \$729 \$1123 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2634 \$1125 \$729 \$451 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2635 b3_r6_b_not \$729 \$291 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2636 \$290 \$729 b3_r6_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2637 \$1201 b3_r6_b \$729 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$2638 \$1200 b3_r6_b_not \$1201 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2639 \$1202 b3_r6_b \$1200 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2640 \$729 b3_r6_b_not \$1202 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2641 \$1203 \$1201 \$1199 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$2642 \$1198 \$1202 \$1203 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2643 \$1204 \$1201 \$1198 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2644 \$1199 \$1202 \$1204 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2645 \$170
+ b2_q0_not|b2_q1_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b4_not|b4_q7_not
+ b4_c7_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2646 \$1129
+ a6_not|b0_p6_not|b1_p6_not|b3_p6_not|b4_p6_not|b5_p6_not|b6_p6_not|b7_p6_not
+ b4_c6_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2647 \$456 a7|b0_p7|b1_p7|b2_p7|b3_p7|b4_p7|b5_p7|b6_p7|b7_p7 \$170 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2648 b4_c7 b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b4|b4_q7 \$456 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2649 \$457 b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b4|b4_q7 b4_c7_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2650 \$172 a7|b0_p7|b1_p7|b2_p7|b3_p7|b4_p7|b5_p7|b6_p7|b7_p7 \$457 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2651 b4_c7
+ b2_q0_not|b2_q1_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b4_not|b4_q7_not
+ \$172 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2652 b4_c6
+ a6_not|b0_p6_not|b1_p6_not|b3_p6_not|b4_p6_not|b5_p6_not|b6_p6_not|b7_p6_not
+ \$1131 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2653 \$224 \$733 \$1129 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2654 \$1131 \$733 \$622 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2655 b4_r6_b_not \$733 \$299 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2656 \$298 \$733 b4_r6_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2657 \$1266 b4_r6_b_not \$1205 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2658 \$733 b4_r6_b_not \$1206 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2659 \$1264 \$1206 \$1207 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2660 \$1265 \$1206 \$1208 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2661 \$177
+ b5_not|b5_q0_not|b5_q1_not|b5_q2_not|b5_q3_not|b5_q4_not|b5_q5_not|b5_q6_not|b5_q7_not
+ b5_c7_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2662 \$1135
+ a6_not|b0_p6_not|b1_p6_not|b3_p6_not|b4_p6_not|b5_p6_not|b6_p6_not|b7_p6_not
+ b5_c6_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2663 \$462 a7|b0_p7|b1_p7|b2_p7|b3_p7|b4_p7|b5_p7|b6_p7|b7_p7 \$177 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2664 b5_c7 b5|b5_q0|b5_q1|b5_q2|b5_q3|b5_q4|b5_q5|b5_q6|b5_q7 \$462 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2665 \$463 b5|b5_q0|b5_q1|b5_q2|b5_q3|b5_q4|b5_q5|b5_q6|b5_q7 b5_c7_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2666 \$179 a7|b0_p7|b1_p7|b2_p7|b3_p7|b4_p7|b5_p7|b6_p7|b7_p7 \$463 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2667 b5_c7
+ b5_not|b5_q0_not|b5_q1_not|b5_q2_not|b5_q3_not|b5_q4_not|b5_q5_not|b5_q6_not|b5_q7_not
+ \$179 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2668 b5_c6
+ a6_not|b0_p6_not|b1_p6_not|b3_p6_not|b4_p6_not|b5_p6_not|b6_p6_not|b7_p6_not
+ \$1137 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2669 \$225 \$737 \$1135 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2670 \$1137 \$737 \$627 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2671 b5_r6_b_not \$737 \$307 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2672 \$306 \$737 b5_r6_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2673 \$1271 b5_r6_b_not \$1209 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2674 \$737 b5_r6_b_not \$1210 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2675 \$1269 \$1210 \$1211 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2676 \$1270 \$1210 \$1212 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2677 \$184
+ b6_not|b6_q0_not|b6_q1_not|b6_q2_not|b6_q3_not|b6_q4_not|b6_q5_not|b6_q6_not|b6_q7_not
+ b6_c7_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2678 \$1141
+ a6_not|b0_p6_not|b1_p6_not|b3_p6_not|b4_p6_not|b5_p6_not|b6_p6_not|b7_p6_not
+ b6_c6_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2679 \$468 a7|b0_p7|b1_p7|b2_p7|b3_p7|b4_p7|b5_p7|b6_p7|b7_p7 \$184 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2680 b6_c7 b6|b6_q0|b6_q1|b6_q2|b6_q3|b6_q4|b6_q5|b6_q6|b6_q7 \$468 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2681 \$469 b6|b6_q0|b6_q1|b6_q2|b6_q3|b6_q4|b6_q5|b6_q6|b6_q7 b6_c7_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2682 \$186 a7|b0_p7|b1_p7|b2_p7|b3_p7|b4_p7|b5_p7|b6_p7|b7_p7 \$469 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2683 b6_c7
+ b6_not|b6_q0_not|b6_q1_not|b6_q2_not|b6_q3_not|b6_q4_not|b6_q5_not|b6_q6_not|b6_q7_not
+ \$186 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2684 b6_c6
+ a6_not|b0_p6_not|b1_p6_not|b3_p6_not|b4_p6_not|b5_p6_not|b6_p6_not|b7_p6_not
+ \$1143 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2685 \$226 \$739 \$1141 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2686 \$1143 \$739 \$632 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2687 b6_r6_b_not \$739 \$315 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2688 \$314 \$739 b6_r6_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2689 \$1276 b6_r6_b_not \$1213 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2690 \$739 b6_r6_b_not \$1214 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2691 \$1274 \$1214 \$1215 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2692 \$1275 \$1214 \$1216 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2693 \$191
+ b7_not|b7_q0_not|b7_q1_not|b7_q2_not|b7_q3_not|b7_q4_not|b7_q5_not|b7_q6_not|b7_q7_not
+ b6_c7_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2694 \$1147
+ a6_not|b0_p6_not|b1_p6_not|b3_p6_not|b4_p6_not|b5_p6_not|b6_p6_not|b7_p6_not
+ b6_c6_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2695 \$474 a7|b0_p7|b1_p7|b2_p7|b3_p7|b4_p7|b5_p7|b6_p7|b7_p7 \$191 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2696 b6_c7 b1_q3|b7|b7_q0|b7_q1|b7_q2|b7_q4|b7_q5|b7_q6|b7_q7 \$474 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2697 \$475 b1_q3|b7|b7_q0|b7_q1|b7_q2|b7_q4|b7_q5|b7_q6|b7_q7 b6_c7_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2698 \$193 a7|b0_p7|b1_p7|b2_p7|b3_p7|b4_p7|b5_p7|b6_p7|b7_p7 \$475 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2699 b6_c7
+ b7_not|b7_q0_not|b7_q1_not|b7_q2_not|b7_q3_not|b7_q4_not|b7_q5_not|b7_q6_not|b7_q7_not
+ \$193 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2700 b6_c6
+ a6_not|b0_p6_not|b1_p6_not|b3_p6_not|b4_p6_not|b5_p6_not|b6_p6_not|b7_p6_not
+ \$1149 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2701 \$227 \$741 \$1147 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2702 \$1149 \$741 \$637 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2703 \$1150 \$741 \$323 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2704 \$322 \$741 \$1151 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2705 \$1281 \$1150 \$1217 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2706 \$741 \$1150 \$1218 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2707 \$1279 \$1218 p13 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2708 \$1280 \$1218 p13_not vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2709 \$1107 \$1110 \$1252 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2710 \$1397 \$1110 \$1253 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2711 \$1403 \$1110 \$1254 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2712 \$1402 \$1110 \$725 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2713 \$1190 b0_r7_b \$725 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$2714 \$1254 b0_r7_b_not \$1190 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2715 \$1191 b0_r7_b \$1254 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2716 \$725 b0_r7_b_not \$1191 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2717 \$1192 \$1190 \$1253 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$2718 \$1252 \$1191 \$1192 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2719 \$1193 \$1190 \$1252 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2720 \$1253 \$1191 \$1193 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2721 \$276 \$1117 \$1257 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2722 \$277 \$1117 \$1258 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2723 \$1412 \$1117 \$1259 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2724 \$1411 \$1117 \$727 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2725 \$1194 b2_r6_b \$727 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$2726 \$1259 b2_r6_b_not \$1194 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2727 \$1195 b2_r6_b \$1259 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2728 \$727 b2_r6_b_not \$1195 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2729 \$1196 \$1194 \$1258 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$2730 \$1257 \$1195 \$1196 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2731 \$1197 \$1194 \$1257 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2732 \$1258 \$1195 \$1197 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2733 \$1198 \$1125 \$285 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2734 \$284 \$1123 \$1198 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2735 \$1199 \$1125 \$284 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2736 \$285 \$1123 \$1199 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2737 \$1200 \$1125 \$1420 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$2738 \$1421 \$1123 \$1200 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2739 \$729 \$1125 \$1421 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2740 \$1420 \$1123 \$729 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2741 \$1264 \$1131 \$293 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2742 \$292 \$1129 \$1264 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2743 \$293 \$1129 \$1265 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2744 \$1266 \$1131 \$1429 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$2745 \$1430 \$1129 \$1266 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2746 \$1429 \$1129 \$733 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2747 \$1205 b4_r6_b \$733 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$2748 \$1206 b4_r6_b \$1266 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2749 \$1207 \$1205 \$1265 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$2750 \$1208 \$1205 \$1264 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2751 \$1269 \$1137 \$301 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2752 \$300 \$1135 \$1269 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2753 \$301 \$1135 \$1270 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2754 \$1271 \$1137 \$1438 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$2755 \$1439 \$1135 \$1271 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2756 \$1438 \$1135 \$737 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2757 \$1209 b5_r6_b \$737 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$2758 \$1210 b5_r6_b \$1271 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2759 \$1211 \$1209 \$1270 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$2760 \$1212 \$1209 \$1269 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2761 \$1274 \$1143 \$309 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2762 \$308 \$1141 \$1274 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2763 \$309 \$1141 \$1275 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2764 \$1276 \$1143 \$1447 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$2765 \$1448 \$1141 \$1276 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2766 \$1447 \$1141 \$739 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2767 \$1213 b6_r6_b \$739 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$2768 \$1214 b6_r6_b \$1276 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2769 \$1215 \$1213 \$1275 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$2770 \$1216 \$1213 \$1274 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2771 \$1279 \$1149 \$317 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2772 \$316 \$1147 \$1279 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2773 \$317 \$1147 \$1280 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2774 \$1281 \$1149 \$1456 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$2775 \$1457 \$1147 \$1281 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2776 \$1456 \$1147 \$741 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2777 \$1217 \$1151 \$741 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2778 \$1218 \$1151 \$1281 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2779 p13 \$1217 \$1280 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2780 p13_not \$1217 \$1279 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2781 \$1397
+ b1_not|b1_q0_not|b1_q1_not|b1_q2_not|b1_q3_not|b1_q4_not|b1_q5_not|b1_q6_not|b1_q7_not
+ b1_c6_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2782 \$1249 a6|b0_p6|b1_p6|b3_p6|b4_p6|b5_p6|b6_p6|b7_p6 \$1397 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2783 b1_c6 b1|b1_q0|b1_q1|b1_q2|b1_q3|b1_q4|b1_q5|b1_q6|b1_q7 \$1249 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2784 \$1250 b1|b1_q0|b1_q1|b1_q2|b1_q3|b1_q4|b1_q5|b1_q6|b1_q7 b1_c6_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2785 \$1107 a6|b0_p6|b1_p6|b3_p6|b4_p6|b5_p6|b6_p6|b7_p6 \$1250 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2786 b1_c6
+ b1_not|b1_q0_not|b1_q1_not|b1_q2_not|b1_q3_not|b1_q4_not|b1_q5_not|b1_q6_not|b1_q7_not
+ \$1107 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2787 \$1110
+ b0_not|b0_q0_not|b0_q1_not|b0_q3_not|b0_q4_not|b0_q5_not|b0_q6_not|b0_q7_not|b1_q2_not
+ b0_c7_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2788 \$1400 a7|b0_p7|b1_p7|b2_p7|b3_p7|b4_p7|b5_p7|b6_p7|b7_p7 \$1110 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2789 b0_c7 b0|b0_q0|b0_q1|b0_q2|b0_q3|b0_q4|b0_q5|b0_q6|b0_q7 \$1400 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2790 \$1401 b0|b0_q0|b0_q1|b0_q2|b0_q3|b0_q4|b0_q5|b0_q6|b0_q7 b0_c7_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2791 \$1112 a7|b0_p7|b1_p7|b2_p7|b3_p7|b4_p7|b5_p7|b6_p7|b7_p7 \$1401 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2792 b0_c7
+ b0_not|b0_q0_not|b0_q1_not|b0_q3_not|b0_q4_not|b0_q5_not|b0_q6_not|b0_q7_not|b1_q2_not
+ \$1112 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2793 \$1252 \$1112 \$1397 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$2794 \$1253 \$1112 \$1107 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2795 \$1254 \$1112 \$1402 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$2796 \$725 \$1112 \$1403 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2797 b0_r7_b_not \$1253 \$275 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2798 \$1255 \$1254 b0_r7_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2799 \$274 \$1252 \$1255 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2800 \$1256 \$1252 \$275 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2801 b0_r7_b \$1254 \$1256 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2802 \$274 \$1253 b0_r7_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2803 \$1117
+ b2_not|b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not
+ b2_c6_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2804 \$1409 a6|b0_p6|b1_p6|b3_p6|b4_p6|b5_p6|b6_p6|b7_p6 \$1117 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2805 b2_c6 b2|b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7 \$1409 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2806 \$1410 b2|b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7 b2_c6_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2807 \$1119 a6|b0_p6|b1_p6|b3_p6|b4_p6|b5_p6|b6_p6|b7_p6 \$1410 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2808 b2_c6
+ b2_not|b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not
+ \$1119 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2809 \$1257 \$1119 \$277 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$2810 \$1258 \$1119 \$276 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2811 \$1259 \$1119 \$1411 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$2812 \$727 \$1119 \$1412 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2813 b2_r6_b_not \$1258 \$283 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2814 \$1260 \$1259 b2_r6_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2815 \$282 \$1257 \$1260 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2816 \$1261 \$1257 \$283 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2817 b2_r6_b \$1259 \$1261 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2818 \$282 \$1258 b2_r6_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2819 \$1123
+ b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b3_not|b3_q0_not|b3_q1_not|b3_q2_not|b3_q3_not|b3_q4_not|b3_q5_not|b3_q6_not|b3_q7_not
+ b3_c6_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2820 \$1418 a6|b0_p6|b1_p6|b3_p6|b4_p6|b5_p6|b6_p6|b7_p6 \$1123 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2821 b3_c6
+ b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b3|b3_q0|b3_q1|b3_q2|b3_q3|b3_q4|b3_q5|b3_q6|b3_q7
+ \$1418 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2822 \$1419
+ b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b3|b3_q0|b3_q1|b3_q2|b3_q3|b3_q4|b3_q5|b3_q6|b3_q7
+ b3_c6_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2823 \$1125 a6|b0_p6|b1_p6|b3_p6|b4_p6|b5_p6|b6_p6|b7_p6 \$1419 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2824 b3_c6
+ b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b3_not|b3_q0_not|b3_q1_not|b3_q2_not|b3_q3_not|b3_q4_not|b3_q5_not|b3_q6_not|b3_q7_not
+ \$1125 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2825 \$223 \$1199 \$1123 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2826 \$1423 \$1200 \$223 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2827 \$1125 \$1198 \$1423 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2828 \$1424 \$1198 \$1123 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2829 \$451 \$1200 \$1424 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2830 \$1125 \$1199 \$451 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2831 b3_r6_b_not \$1199 \$291 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2832 \$1262 \$1200 b3_r6_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2833 \$290 \$1198 \$1262 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2834 \$1263 \$1198 \$291 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2835 b3_r6_b \$1200 \$1263 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2836 \$290 \$1199 b3_r6_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2837 \$1265 \$1131 \$292 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2838 \$733 \$1131 \$1430 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2839 \$224 \$1265 \$1129 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2840 \$1432 \$1266 \$224 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2841 \$1131 \$1264 \$1432 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2842 \$1433 \$1264 \$1129 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2843 \$622 \$1266 \$1433 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2844 \$1131 \$1265 \$622 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2845 b4_r6_b_not \$1265 \$299 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2846 \$1267 \$1266 b4_r6_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2847 \$298 \$1264 \$1267 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2848 \$1268 \$1264 \$299 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2849 b4_r6_b \$1266 \$1268 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2850 \$298 \$1265 b4_r6_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2851 \$1270 \$1137 \$300 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2852 \$737 \$1137 \$1439 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2853 \$225 \$1270 \$1135 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2854 \$1441 \$1271 \$225 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2855 \$1137 \$1269 \$1441 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2856 \$1442 \$1269 \$1135 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2857 \$627 \$1271 \$1442 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2858 \$1137 \$1270 \$627 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2859 b5_r6_b_not \$1270 \$307 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2860 \$1272 \$1271 b5_r6_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2861 \$306 \$1269 \$1272 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2862 \$1273 \$1269 \$307 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2863 b5_r6_b \$1271 \$1273 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2864 \$306 \$1270 b5_r6_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2865 \$1141
+ b6_not|b6_q0_not|b6_q1_not|b6_q2_not|b6_q3_not|b6_q4_not|b6_q5_not|b6_q6_not|b6_q7_not
+ b6_c6_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2866 \$1445 a6|b0_p6|b1_p6|b3_p6|b4_p6|b5_p6|b6_p6|b7_p6 \$1141 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2867 b6_c6 b6|b6_q0|b6_q1|b6_q2|b6_q3|b6_q4|b6_q5|b6_q6|b6_q7 \$1445 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2868 \$1446 b6|b6_q0|b6_q1|b6_q2|b6_q3|b6_q4|b6_q5|b6_q6|b6_q7 b6_c6_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2869 \$1143 a6|b0_p6|b1_p6|b3_p6|b4_p6|b5_p6|b6_p6|b7_p6 \$1446 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2870 b6_c6
+ b6_not|b6_q0_not|b6_q1_not|b6_q2_not|b6_q3_not|b6_q4_not|b6_q5_not|b6_q6_not|b6_q7_not
+ \$1143 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2871 \$1275 \$1143 \$308 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2872 \$739 \$1143 \$1448 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2873 \$226 \$1275 \$1141 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2874 \$1450 \$1276 \$226 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2875 \$1143 \$1274 \$1450 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2876 \$1451 \$1274 \$1141 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2877 \$632 \$1276 \$1451 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2878 \$1143 \$1275 \$632 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2879 b6_r6_b_not \$1275 \$315 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2880 \$1277 \$1276 b6_r6_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2881 \$314 \$1274 \$1277 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2882 \$1278 \$1274 \$315 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2883 b6_r6_b \$1276 \$1278 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2884 \$314 \$1275 b6_r6_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2885 \$1147
+ b7_not|b7_q0_not|b7_q1_not|b7_q2_not|b7_q3_not|b7_q4_not|b7_q5_not|b7_q6_not|b7_q7_not
+ b6_c6_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2886 \$1454 a6|b0_p6|b1_p6|b3_p6|b4_p6|b5_p6|b6_p6|b7_p6 \$1147 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2887 b6_c6 b1_q3|b7|b7_q0|b7_q1|b7_q2|b7_q4|b7_q5|b7_q6|b7_q7 \$1454 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2888 \$1455 b1_q3|b7|b7_q0|b7_q1|b7_q2|b7_q4|b7_q5|b7_q6|b7_q7 b6_c6_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2889 \$1149 a6|b0_p6|b1_p6|b3_p6|b4_p6|b5_p6|b6_p6|b7_p6 \$1455 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2890 b6_c6
+ b7_not|b7_q0_not|b7_q1_not|b7_q2_not|b7_q3_not|b7_q4_not|b7_q5_not|b7_q6_not|b7_q7_not
+ \$1149 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2891 \$1280 \$1149 \$316 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2892 \$741 \$1149 \$1457 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2893 \$227 \$1280 \$1147 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2894 \$1459 \$1281 \$227 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2895 \$1149 \$1279 \$1459 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2896 \$1460 \$1279 \$1147 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2897 \$637 \$1281 \$1460 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2898 \$1149 \$1280 \$637 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2899 \$1150 \$1280 \$323 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2900 \$1282 \$1281 \$1150 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2901 \$322 \$1279 \$1282 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2902 \$1283 \$1279 \$323 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2903 \$1151 \$1281 \$1283 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2904 \$322 \$1280 \$1151 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2905 \$2358
+ a5_not|b0_p5_not|b1_p5_not|b2_p5_not|b3_p5_not|b5_p5_not|b6_p5_not|b7_p5_not
+ b1_c5_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2906 b1_c5
+ a5_not|b0_p5_not|b1_p5_not|b2_p5_not|b3_p5_not|b5_p5_not|b6_p5_not|b7_p5_not
+ \$2083 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2907 \$2085
+ a6_not|b0_p6_not|b1_p6_not|b3_p6_not|b4_p6_not|b5_p6_not|b6_p6_not|b7_p6_not
+ b0_c6_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2908 b0_c6
+ a6_not|b0_p6_not|b1_p6_not|b3_p6_not|b4_p6_not|b5_p6_not|b6_p6_not|b7_p6_not
+ \$2086 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2909 \$2083 \$2085 \$2208 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2910 \$2358 \$2085 \$2210 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2911 \$2361 \$2085 \$2209 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2912 \$2360 \$2085 \$2068 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2913 \$221 \$1253 \$1110 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2914 \$1402 \$2068 \$2085 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2915 \$1405 \$1254 \$221 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2916 \$1112 \$1252 \$1405 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2917 \$1406 \$1252 \$1110 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2918 \$608 \$1254 \$1406 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2919 \$1112 \$1253 \$608 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2920 \$2086 \$2068 \$1403 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2921 b0_r6_b_not \$2068 \$1191 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2922 \$1190 \$2068 b0_r6_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2923 \$2090
+ a5_not|b0_p5_not|b1_p5_not|b2_p5_not|b3_p5_not|b5_p5_not|b6_p5_not|b7_p5_not
+ b2_c5_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2924 b2_c5
+ a5_not|b0_p5_not|b1_p5_not|b2_p5_not|b3_p5_not|b5_p5_not|b6_p5_not|b7_p5_not
+ \$2091 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2925 \$1192 \$2090 \$2215 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2926 \$1193 \$2090 \$2217 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2927 \$2369 \$2090 \$2216 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2928 \$2368 \$2090 \$2070 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2929 \$222 \$1258 \$1117 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2930 \$1411 \$2070 \$2090 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2931 \$1414 \$1259 \$222 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2932 \$1119 \$1257 \$1414 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2933 \$1415 \$1257 \$1117 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2934 \$613 \$1259 \$1415 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2935 \$1119 \$1258 \$613 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2936 \$2091 \$2070 \$1412 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2937 b2_r5_b_not \$2070 \$1195 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2938 \$1194 \$2070 b2_r5_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2939 \$2095
+ a5_not|b0_p5_not|b1_p5_not|b2_p5_not|b3_p5_not|b5_p5_not|b6_p5_not|b7_p5_not
+ b2_c5_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2940 b3_c5
+ a5_not|b0_p5_not|b1_p5_not|b2_p5_not|b3_p5_not|b5_p5_not|b6_p5_not|b7_p5_not
+ \$2096 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2941 \$2162 \$2096 \$1197 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$2942 \$1196 \$2095 \$2162 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2943 \$2163 \$2096 \$1196 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2944 \$1197 \$2095 \$2163 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2945 \$2164 \$2096 \$2375 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$2946 \$2376 \$2095 \$2164 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2947 \$2072 \$2096 \$2376 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2948 \$2375 \$2095 \$2072 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2949 \$1420 \$2072 \$2095 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2950 \$2096 \$2072 \$1421 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2951 b3_r5_b_not \$2072 \$1202 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2952 \$1201 \$2072 b3_r5_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2953 \$2165 b3_r5_b \$2072 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$2954 \$2164 b3_r5_b_not \$2165 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2955 \$2166 b3_r5_b \$2164 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2956 \$2072 b3_r5_b_not \$2166 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2957 \$2167 \$2165 \$2163 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$2958 \$2162 \$2166 \$2167 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2959 \$2168 \$2165 \$2162 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$2960 \$2163 \$2166 \$2168 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2961 \$2100
+ a5_not|b0_p5_not|b1_p5_not|b2_p5_not|b3_p5_not|b5_p5_not|b6_p5_not|b7_p5_not
+ b2_c5_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2962 \$1129
+ b2_q0_not|b2_q1_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b4_not|b4_q7_not
+ b4_c6_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2963 \$1427 a6|b0_p6|b1_p6|b3_p6|b4_p6|b5_p6|b6_p6|b7_p6 \$1129 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2964 b4_c6 b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b4|b4_q7 \$1427 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2965 \$1428 b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b4|b4_q7 b4_c6_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2966 \$1131 a6|b0_p6|b1_p6|b3_p6|b4_p6|b5_p6|b6_p6|b7_p6 \$1428 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2967 \$2102
+ a5_not|b0_p5_not|b1_p5_not|b2_p5_not|b3_p5_not|b5_p5_not|b6_p5_not|b7_p5_not
+ \$2101 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2968 b4_c6
+ b2_q0_not|b2_q1_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b4_not|b4_q7_not
+ \$1131 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2969 \$1203 \$2100 \$2169 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2970 \$1204 \$2100 \$2224 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2971 \$2384 \$2100 \$2170 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2972 \$2383 \$2100 \$2074 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2973 \$1429 \$2074 \$2100 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2974 \$2101 \$2074 \$1430 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2975 b4_r5_b_not \$2074 \$1206 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2976 \$1205 \$2074 b4_r5_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2977 \$2170 b4_r5_b_not \$2225 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2978 \$2169 \$2226 \$2227 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2979 \$2106
+ a5_not|b0_p5_not|b1_p5_not|b2_p5_not|b3_p5_not|b5_p5_not|b6_p5_not|b7_p5_not
+ \$2105 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2980 \$1135
+ b5_not|b5_q0_not|b5_q1_not|b5_q2_not|b5_q3_not|b5_q4_not|b5_q5_not|b5_q6_not|b5_q7_not
+ b5_c6_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2981 \$1436 a6|b0_p6|b1_p6|b3_p6|b4_p6|b5_p6|b6_p6|b7_p6 \$1135 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2982 b5_c6 b5|b5_q0|b5_q1|b5_q2|b5_q3|b5_q4|b5_q5|b5_q6|b5_q7 \$1436 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2983 \$1437 b5|b5_q0|b5_q1|b5_q2|b5_q3|b5_q4|b5_q5|b5_q6|b5_q7 b5_c6_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2984 \$1137 a6|b0_p6|b1_p6|b3_p6|b4_p6|b5_p6|b6_p6|b7_p6 \$1437 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2985 b5_c5
+ a5_not|b0_p5_not|b1_p5_not|b2_p5_not|b3_p5_not|b5_p5_not|b6_p5_not|b7_p5_not
+ \$2107 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2986 b5_c6
+ b5_not|b5_q0_not|b5_q1_not|b5_q2_not|b5_q3_not|b5_q4_not|b5_q5_not|b5_q6_not|b5_q7_not
+ \$1137 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2987 \$1207 \$2106 \$2171 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2988 \$1208 \$2106 \$2229 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2989 \$2392 \$2106 \$2172 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2990 \$2391 \$2106 \$2076 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$2991 \$1438 \$2076 \$2106 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2992 \$2107 \$2076 \$1439 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$2993 b5_r5_b_not \$2076 \$1210 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2994 \$1209 \$2076 b5_r5_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$2995 \$2172 b5_r5_b_not \$2230 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2996 \$2171 \$2231 \$2232 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$2997 \$2111
+ a5_not|b0_p5_not|b1_p5_not|b2_p5_not|b3_p5_not|b5_p5_not|b6_p5_not|b7_p5_not
+ b6_c5_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$2998 b6_c5
+ a5_not|b0_p5_not|b1_p5_not|b2_p5_not|b3_p5_not|b5_p5_not|b6_p5_not|b7_p5_not
+ \$2112 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$2999 \$1211 \$2111 \$2173 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3000 \$1212 \$2111 \$2236 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3001 \$2399 \$2111 \$2174 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3002 \$2398 \$2111 \$2078 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3003 \$1447 \$2078 \$2111 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3004 \$2112 \$2078 \$1448 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3005 b6_r5_b_not \$2078 \$1214 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3006 \$1213 \$2078 b6_r5_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3007 \$2174 b6_r5_b_not \$2237 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3008 \$2173 \$2238 \$2239 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3009 \$2116
+ a5_not|b0_p5_not|b1_p5_not|b2_p5_not|b3_p5_not|b5_p5_not|b6_p5_not|b7_p5_not
+ \$2115 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3010 b6_c5
+ a5_not|b0_p5_not|b1_p5_not|b2_p5_not|b3_p5_not|b5_p5_not|b6_p5_not|b7_p5_not
+ \$2117 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3011 \$1215 \$2116 \$2175 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3012 \$1216 \$2116 \$2241 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3013 \$2407 \$2116 \$2176 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3014 \$2406 \$2116 \$2080 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3015 \$1456 \$2080 \$2116 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3016 \$2117 \$2080 \$1457 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3017 \$2118 \$2080 \$1218 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3018 \$1217 \$2080 \$2119 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3019 \$2176 \$2118 \$2242 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3020 \$2175 \$2243 p12 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3021 \$2358
+ b1_not|b1_q0_not|b1_q1_not|b1_q2_not|b1_q3_not|b1_q4_not|b1_q5_not|b1_q6_not|b1_q7_not
+ b1_c5_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3022 \$2202 a5|b0_p5|b1_p5|b3_p5|b4_p5|b5_p5|b6_p5|b7_p5 \$2358 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3023 b1_c5 b1|b1_q0|b1_q1|b1_q2|b1_q3|b1_q4|b1_q5|b1_q6|b1_q7 \$2202 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3024 \$2204 b1|b1_q0|b1_q1|b1_q2|b1_q3|b1_q4|b1_q5|b1_q6|b1_q7 b1_c5_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3025 \$2083 a5|b0_p5|b1_p5|b3_p5|b4_p5|b5_p5|b6_p5|b7_p5 \$2204 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3026 b1_c5
+ b1_not|b1_q0_not|b1_q1_not|b1_q2_not|b1_q3_not|b1_q4_not|b1_q5_not|b1_q6_not|b1_q7_not
+ \$2083 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3027 \$2208 \$2086 \$2358 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3028 \$2210 \$2086 \$2083 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3029 \$2209 \$2086 \$2360 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3030 \$2068 \$2086 \$2361 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3031 \$2211 b0_r6_b \$2068 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3032 \$2209 b0_r6_b_not \$2211 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3033 \$2212 b0_r6_b \$2209 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3034 \$2068 b0_r6_b_not \$2212 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3035 \$2213 \$2211 \$2210 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3036 \$2208 \$2212 \$2213 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3037 \$2214 \$2211 \$2208 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3038 \$2210 \$2212 \$2214 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3039 \$2215 \$2091 \$1193 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3040 \$2217 \$2091 \$1192 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3041 \$2216 \$2091 \$2368 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3042 \$2070 \$2091 \$2369 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3043 \$2218 b2_r5_b \$2070 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3044 \$2216 b2_r5_b_not \$2218 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3045 \$2219 b2_r5_b \$2216 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3046 \$2070 b2_r5_b_not \$2219 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3047 \$2220 \$2218 \$2217 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3048 \$2215 \$2219 \$2220 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3049 \$2221 \$2218 \$2215 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3050 \$2217 \$2219 \$2221 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3051 \$2095
+ b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b3_not|b3_q0_not|b3_q1_not|b3_q2_not|b3_q3_not|b3_q4_not|b3_q5_not|b3_q6_not|b3_q7_not
+ b2_c5_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3052 \$2222 a5|b0_p5|b1_p5|b3_p5|b4_p5|b5_p5|b6_p5|b7_p5 \$2095 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3053 b3_c5
+ b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b3|b3_q0|b3_q1|b3_q2|b3_q3|b3_q4|b3_q5|b3_q6|b3_q7
+ \$2222 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3054 \$2223
+ b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b3|b3_q0|b3_q1|b3_q2|b3_q3|b3_q4|b3_q5|b3_q6|b3_q7
+ b2_c5_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3055 \$2096 a5|b0_p5|b1_p5|b3_p5|b4_p5|b5_p5|b6_p5|b7_p5 \$2223 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3056 b3_c5
+ b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b3_not|b3_q0_not|b3_q1_not|b3_q2_not|b3_q3_not|b3_q4_not|b3_q5_not|b3_q6_not|b3_q7_not
+ \$2096 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3057 \$2169 \$2101 \$1204 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3058 \$2224 \$2101 \$1203 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3059 \$2170 \$2101 \$2383 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3060 \$2074 \$2101 \$2384 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3061 \$2225 b4_r5_b \$2074 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3062 \$2226 b4_r5_b \$2170 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3063 \$2074 b4_r5_b_not \$2226 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3064 \$2227 \$2225 \$2224 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3065 \$2228 \$2225 \$2169 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3066 \$2224 \$2226 \$2228 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3067 \$2171 \$2107 \$1208 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3068 \$2229 \$2107 \$1207 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3069 \$2172 \$2107 \$2391 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3070 \$2076 \$2107 \$2392 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3071 \$2230 b5_r5_b \$2076 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3072 \$2231 b5_r5_b \$2172 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3073 \$2076 b5_r5_b_not \$2231 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3074 \$2232 \$2230 \$2229 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3075 \$2233 \$2230 \$2171 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3076 \$2229 \$2231 \$2233 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3077 \$2173 \$2112 \$1212 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3078 \$2236 \$2112 \$1211 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3079 \$2174 \$2112 \$2398 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3080 \$2078 \$2112 \$2399 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3081 \$2237 b6_r5_b \$2078 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3082 \$2238 b6_r5_b \$2174 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3083 \$2078 b6_r5_b_not \$2238 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3084 \$2239 \$2237 \$2236 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3085 \$2240 \$2237 \$2173 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3086 \$2236 \$2238 \$2240 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3087 \$2175 \$2117 \$1216 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3088 \$2241 \$2117 \$1215 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3089 \$2176 \$2117 \$2406 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3090 \$2080 \$2117 \$2407 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3091 \$2242 \$2119 \$2080 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3092 \$2243 \$2119 \$2176 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3093 \$2080 \$2118 \$2243 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3094 p12 \$2242 \$2241 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$3095 p12_not \$2242 \$2175 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3096 \$2241 \$2243 p12_not vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3097 \$2085
+ b0_not|b0_q0_not|b0_q1_not|b0_q3_not|b0_q4_not|b0_q5_not|b0_q6_not|b0_q7_not|b1_q2_not
+ b0_c6_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3098 \$2205 a6|b0_p6|b1_p6|b3_p6|b4_p6|b5_p6|b6_p6|b7_p6 \$2085 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3099 b0_c6 b0|b0_q0|b0_q1|b0_q2|b0_q3|b0_q4|b0_q5|b0_q6|b0_q7 \$2205 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3100 \$2207 b0|b0_q0|b0_q1|b0_q2|b0_q3|b0_q4|b0_q5|b0_q6|b0_q7 b0_c6_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3101 \$2086 a6|b0_p6|b1_p6|b3_p6|b4_p6|b5_p6|b6_p6|b7_p6 \$2207 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3102 b0_c6
+ b0_not|b0_q0_not|b0_q1_not|b0_q3_not|b0_q4_not|b0_q5_not|b0_q6_not|b0_q7_not|b1_q2_not
+ \$2086 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3103 \$2111
+ b6_not|b6_q0_not|b6_q1_not|b6_q2_not|b6_q3_not|b6_q4_not|b6_q5_not|b6_q6_not|b6_q7_not
+ b6_c5_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3104 \$2234 a5|b0_p5|b1_p5|b3_p5|b4_p5|b5_p5|b6_p5|b7_p5 \$2111 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3105 b6_c5 b6|b6_q0|b6_q1|b6_q2|b6_q3|b6_q4|b6_q5|b6_q6|b6_q7 \$2234 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3106 \$2235 b6|b6_q0|b6_q1|b6_q2|b6_q3|b6_q4|b6_q5|b6_q6|b6_q7 b6_c5_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3107 \$2112 a5|b0_p5|b1_p5|b3_p5|b4_p5|b5_p5|b6_p5|b7_p5 \$2235 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3108 b6_c5
+ b6_not|b6_q0_not|b6_q1_not|b6_q2_not|b6_q3_not|b6_q4_not|b6_q5_not|b6_q6_not|b6_q7_not
+ \$2112 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3109 \$2090
+ b2_not|b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not
+ b2_c5_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3110 \$2366 a5|b0_p5|b1_p5|b3_p5|b4_p5|b5_p5|b6_p5|b7_p5 \$2090 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3111 b2_c5 b2|b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7 \$2366 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3112 \$2367 b2|b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7 b2_c5_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3113 \$2091 a5|b0_p5|b1_p5|b3_p5|b4_p5|b5_p5|b6_p5|b7_p5 \$2367 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3114 b2_c5
+ b2_not|b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not
+ \$2091 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3115 \$2100
+ b2_q0_not|b2_q1_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b4_not|b4_q7_not
+ b2_c5_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3116 \$2381 a5|b0_p5|b1_p5|b3_p5|b4_p5|b5_p5|b6_p5|b7_p5 \$2100 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3117 \$2102 b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b4|b4_q7 \$2381 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3118 \$2382 b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b4|b4_q7 b2_c5_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3119 \$2101 a5|b0_p5|b1_p5|b3_p5|b4_p5|b5_p5|b6_p5|b7_p5 \$2382 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3120 \$2102
+ b2_q0_not|b2_q1_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b4_not|b4_q7_not
+ \$2101 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3121 \$2106
+ b5_not|b5_q0_not|b5_q1_not|b5_q2_not|b5_q3_not|b5_q4_not|b5_q5_not|b5_q6_not|b5_q7_not
+ \$2105 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3122 \$2389 a5|b0_p5|b1_p5|b3_p5|b4_p5|b5_p5|b6_p5|b7_p5 \$2106 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3123 b5_c5 b5|b5_q0|b5_q1|b5_q2|b5_q3|b5_q4|b5_q5|b5_q6|b5_q7 \$2389 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3124 \$2390 b5|b5_q0|b5_q1|b5_q2|b5_q3|b5_q4|b5_q5|b5_q6|b5_q7 \$2105 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3125 \$2107 a5|b0_p5|b1_p5|b3_p5|b4_p5|b5_p5|b6_p5|b7_p5 \$2390 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3126 b5_c5
+ b5_not|b5_q0_not|b5_q1_not|b5_q2_not|b5_q3_not|b5_q4_not|b5_q5_not|b5_q6_not|b5_q7_not
+ \$2107 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3127 \$2116
+ b7_not|b7_q0_not|b7_q1_not|b7_q2_not|b7_q3_not|b7_q4_not|b7_q5_not|b7_q6_not|b7_q7_not
+ \$2115 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3128 \$2404 a5|b0_p5|b1_p5|b3_p5|b4_p5|b5_p5|b6_p5|b7_p5 \$2116 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3129 b6_c5 b1_q3|b7|b7_q0|b7_q1|b7_q2|b7_q4|b7_q5|b7_q6|b7_q7 \$2404 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3130 \$2405 b1_q3|b7|b7_q0|b7_q1|b7_q2|b7_q4|b7_q5|b7_q6|b7_q7 \$2115 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3131 \$2117 a5|b0_p5|b1_p5|b3_p5|b4_p5|b5_p5|b6_p5|b7_p5 \$2405 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3132 b6_c5
+ b7_not|b7_q0_not|b7_q1_not|b7_q2_not|b7_q3_not|b7_q4_not|b7_q5_not|b7_q6_not|b7_q7_not
+ \$2117 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3133 \$1402 \$2210 \$2085 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3134 \$2362 \$2209 \$1402 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3135 \$2086 \$2208 \$2362 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3136 \$2363 \$2208 \$2085 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3137 \$1403 \$2209 \$2363 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3138 \$2086 \$2210 \$1403 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3139 \$1411 \$2217 \$2090 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3140 \$2370 \$2216 \$1411 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3141 \$2091 \$2215 \$2370 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3142 \$2371 \$2215 \$2090 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3143 \$1412 \$2216 \$2371 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3144 \$2091 \$2217 \$1412 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3145 \$1420 \$2163 \$2095 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3146 \$2377 \$2164 \$1420 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3147 \$2096 \$2162 \$2377 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3148 \$2378 \$2162 \$2095 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3149 \$1421 \$2164 \$2378 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3150 \$2096 \$2163 \$1421 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3151 b3_r5_b_not \$2163 \$1202 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3152 \$2379 \$2164 b3_r5_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3153 \$1201 \$2162 \$2379 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3154 \$2380 \$2162 \$1202 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3155 b3_r5_b \$2164 \$2380 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3156 \$1201 \$2163 b3_r5_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3157 \$1429 \$2224 \$2100 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3158 \$2385 \$2170 \$1429 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3159 \$2101 \$2169 \$2385 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3160 \$2386 \$2169 \$2100 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3161 \$1430 \$2170 \$2386 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3162 \$2101 \$2224 \$1430 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3163 \$1438 \$2229 \$2106 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3164 \$2393 \$2172 \$1438 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3165 \$2107 \$2171 \$2393 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3166 \$2394 \$2171 \$2106 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3167 \$1439 \$2172 \$2394 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3168 \$2107 \$2229 \$1439 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3169 \$1447 \$2236 \$2111 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3170 \$2400 \$2174 \$1447 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3171 \$2112 \$2173 \$2400 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3172 \$2401 \$2173 \$2111 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3173 \$1448 \$2174 \$2401 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3174 \$2112 \$2236 \$1448 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3175 \$1456 \$2241 \$2116 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3176 \$2408 \$2176 \$1456 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3177 \$2117 \$2175 \$2408 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3178 \$2409 \$2175 \$2116 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3179 \$1457 \$2176 \$2409 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3180 \$2117 \$2241 \$1457 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3181 \$3115
+ a4_not|b0_p4_not|b1_p4_not|b2_p4_not|b3_p4_not|b5_p4_not|b6_p4_not|b7_p4_not
+ b1_c4_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3182 b1_c4
+ a4_not|b0_p4_not|b1_p4_not|b2_p4_not|b3_p4_not|b5_p4_not|b6_p4_not|b7_p4_not
+ \$3043 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3183 \$3045
+ a5_not|b0_p5_not|b1_p5_not|b2_p5_not|b3_p5_not|b5_p5_not|b6_p5_not|b7_p5_not
+ b0_c5_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3184 b0_c5
+ a5_not|b0_p5_not|b1_p5_not|b2_p5_not|b3_p5_not|b5_p5_not|b6_p5_not|b7_p5_not
+ \$3047 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3185 \$2360 \$3034 \$3045 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3186 \$3047 \$3034 \$2361 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3187 b0_r5_b_not \$3034 \$2212 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3188 b0_r6_b_not \$2210 \$1191 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3189 \$2364 \$2209 b0_r6_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3190 \$1190 \$2208 \$2364 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3191 \$2365 \$2208 \$1191 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3192 b0_r6_b \$2209 \$2365 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3193 \$2211 \$3034 b0_r5_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3194 \$1190 \$2210 b0_r6_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3195 \$3051
+ a4_not|b0_p4_not|b1_p4_not|b2_p4_not|b3_p4_not|b5_p4_not|b6_p4_not|b7_p4_not
+ b2_c4_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3196 b2_c4
+ a4_not|b0_p4_not|b1_p4_not|b2_p4_not|b3_p4_not|b5_p4_not|b6_p4_not|b7_p4_not
+ \$3053 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3197 \$2368 \$3035 \$3051 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3198 \$3053 \$3035 \$2369 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3199 b2_r4_b_not \$3035 \$2219 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3200 b2_r5_b_not \$2217 \$1195 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3201 \$2372 \$2216 b2_r5_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3202 \$1194 \$2215 \$2372 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3203 \$2373 \$2215 \$1195 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3204 b2_r5_b \$2216 \$2373 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3205 \$2218 \$3035 b2_r4_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3206 \$1194 \$2217 b2_r5_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3207 \$3057
+ a4_not|b0_p4_not|b1_p4_not|b2_p4_not|b3_p4_not|b5_p4_not|b6_p4_not|b7_p4_not
+ b2_c4_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3208 b2_c4
+ a4_not|b0_p4_not|b1_p4_not|b2_p4_not|b3_p4_not|b5_p4_not|b6_p4_not|b7_p4_not
+ \$3058 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3209 \$2220 \$3057 \$3189 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3210 \$2221 \$3057 \$3191 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3211 \$3342 \$3057 \$3190 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3212 \$3118 \$3057 \$3036 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3213 \$2375 \$3036 \$3057 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3214 \$3058 \$3036 \$2376 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3215 b3_r4_b_not \$3036 \$2166 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3216 \$2165 \$3036 b3_r4_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3217 \$3119 b3_r4_b \$3036 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3218 \$3190 b3_r4_b_not \$3119 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3219 \$3120 b3_r4_b \$3190 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3220 \$3036 b3_r4_b_not \$3120 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3221 \$3121 \$3119 \$3191 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3222 \$3189 \$3120 \$3121 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3223 \$3122 \$3119 \$3189 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3224 \$3191 \$3120 \$3122 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3225 \$3062
+ a4_not|b0_p4_not|b1_p4_not|b2_p4_not|b3_p4_not|b5_p4_not|b6_p4_not|b7_p4_not
+ b2_c4_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3226 b2_c4
+ a4_not|b0_p4_not|b1_p4_not|b2_p4_not|b3_p4_not|b5_p4_not|b6_p4_not|b7_p4_not
+ \$3064 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3227 \$2383 \$3037 \$3062 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3228 \$3064 \$3037 \$2384 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3229 b4_r4_b_not \$3037 \$2226 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3230 b4_r5_b_not \$2224 \$1206 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3231 \$2387 \$2170 b4_r5_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3232 \$1205 \$2169 \$2387 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3233 \$2388 \$2169 \$1206 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3234 b4_r5_b \$2170 \$2388 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3235 \$2225 \$3037 b4_r4_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3236 \$1205 \$2224 b4_r5_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3237 \$3193 b4_r4_b_not \$3195 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3238 \$3192 \$3124 \$3196 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3239 \$3068
+ a4_not|b0_p4_not|b1_p4_not|b2_p4_not|b3_p4_not|b5_p4_not|b6_p4_not|b7_p4_not
+ \$3067 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3240 \$3071
+ a4_not|b0_p4_not|b1_p4_not|b2_p4_not|b3_p4_not|b5_p4_not|b6_p4_not|b7_p4_not
+ \$3070 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3241 \$2391 \$3038 \$3068 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3242 \$3070 \$3038 \$2392 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3243 b5_r4_b_not \$3038 \$2231 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3244 b5_r5_b_not \$2229 \$1210 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3245 \$2395 \$2172 b5_r5_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3246 \$1209 \$2171 \$2395 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3247 \$2396 \$2171 \$1210 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3248 b5_r5_b \$2172 \$2396 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3249 \$2230 \$3038 b5_r4_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3250 \$1209 \$2229 b5_r5_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3251 \$3198 b5_r4_b_not \$3200 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3252 \$3197 \$3127 \$3201 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3253 \$3075
+ a4_not|b0_p4_not|b1_p4_not|b2_p4_not|b3_p4_not|b5_p4_not|b6_p4_not|b7_p4_not
+ b6_c4_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3254 b6_c4
+ a4_not|b0_p4_not|b1_p4_not|b2_p4_not|b3_p4_not|b5_p4_not|b6_p4_not|b7_p4_not
+ \$3077 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3255 \$2398 \$3039 \$3075 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3256 \$3077 \$3039 \$2399 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3257 b6_r4_b_not \$3039 \$2238 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3258 b6_r5_b_not \$2236 \$1214 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3259 \$2402 \$2174 b6_r5_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3260 \$1213 \$2173 \$2402 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3261 \$2403 \$2173 \$1214 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3262 b6_r5_b \$2174 \$2403 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3263 \$2237 \$3039 b6_r4_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3264 \$1213 \$2236 b6_r5_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3265 \$3203 b6_r4_b_not \$3205 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3266 \$3202 \$3130 \$3206 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3267 \$3081
+ a4_not|b0_p4_not|b1_p4_not|b2_p4_not|b3_p4_not|b5_p4_not|b6_p4_not|b7_p4_not
+ \$3080 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3268 \$3084
+ a4_not|b0_p4_not|b1_p4_not|b2_p4_not|b3_p4_not|b5_p4_not|b6_p4_not|b7_p4_not
+ \$3083 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3269 \$2406 \$3040 \$3081 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3270 \$3083 \$3040 \$2407 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3271 \$3085 \$3040 \$2243 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3272 \$2118 \$2241 \$1218 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3273 \$2410 \$2176 \$2118 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3274 \$1217 \$2175 \$2410 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3275 \$2411 \$2175 \$1218 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3276 \$2119 \$2176 \$2411 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3277 \$2242 \$3040 \$3086 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3278 \$1217 \$2241 \$2119 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3279 \$3208 \$3085 \$3210 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3280 \$3207 \$3133 p11 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3281 \$3043 \$3045 \$3175 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3282 \$3328 \$3045 \$3176 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3283 \$3178 b0_r5_b \$3034 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3284 \$3176 b0_r5_b_not \$3178 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3285 \$3034 b0_r5_b_not \$3179 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3286 \$3180 \$3178 \$3177 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3287 \$3175 \$3179 \$3180 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3288 \$3177 \$3179 \$3181 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3289 \$2213 \$3051 \$3182 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3290 \$3335 \$3051 \$3183 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3291 \$3185 b2_r4_b \$3035 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3292 \$3183 b2_r4_b_not \$3185 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3293 \$3035 b2_r4_b_not \$3186 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3294 \$3187 \$3185 \$3184 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3295 \$3182 \$3186 \$3187 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3296 \$3184 \$3186 \$3188 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3297 \$3189 \$3058 \$2221 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3298 \$3191 \$3058 \$2220 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3299 \$3190 \$3058 \$3118 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3300 \$3036 \$3058 \$3342 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3301 \$2167 \$3062 \$3192 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3302 \$2168 \$3062 \$3194 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3303 \$3349 \$3062 \$3193 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3304 \$3123 \$3062 \$3037 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3305 \$3195 b4_r4_b \$3037 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3306 \$3124 b4_r4_b \$3193 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3307 \$3037 b4_r4_b_not \$3124 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3308 \$3196 \$3195 \$3194 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3309 \$3125 \$3195 \$3192 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3310 \$3194 \$3124 \$3125 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3311 \$2227 \$3068 \$3197 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3312 \$2228 \$3068 \$3199 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3313 \$3356 \$3068 \$3198 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3314 \$3126 \$3068 \$3038 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3315 \$3200 b5_r4_b \$3038 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3316 \$3127 b5_r4_b \$3198 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3317 \$3038 b5_r4_b_not \$3127 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3318 \$3201 \$3200 \$3199 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3319 \$3128 \$3200 \$3197 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3320 \$3199 \$3127 \$3128 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3321 \$2232 \$3075 \$3202 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3322 \$2233 \$3075 \$3204 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3323 \$3364 \$3075 \$3203 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3324 \$3129 \$3075 \$3039 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3325 \$3205 b6_r4_b \$3039 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3326 \$3130 b6_r4_b \$3203 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3327 \$3039 b6_r4_b_not \$3130 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3328 \$3206 \$3205 \$3204 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3329 \$3131 \$3205 \$3202 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3330 \$3204 \$3130 \$3131 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3331 \$2239 \$3081 \$3207 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3332 \$2240 \$3081 \$3209 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3333 \$3371 \$3081 \$3208 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3334 \$3132 \$3081 \$3040 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3335 \$3210 \$3086 \$3040 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3336 \$3133 \$3086 \$3208 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3337 \$3040 \$3085 \$3133 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3338 p11 \$3210 \$3209 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$3339 p11_not \$3210 \$3207 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3340 \$3209 \$3133 p11_not vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3341 \$3115
+ b1_not|b1_q0_not|b1_q1_not|b1_q2_not|b1_q3_not|b1_q4_not|b1_q5_not|b1_q6_not|b1_q7_not
+ b1_c4_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3342 \$3323 a4|b0_p4|b1_p4|b2_p4|b3_p4|b4_p4|b5_p4|b6_p4|b7_p4 \$3115 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3343 b1_c4 b1|b1_q0|b1_q1|b1_q2|b1_q3|b1_q4|b1_q5|b1_q6|b1_q7 \$3323 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3344 \$3324 b1|b1_q0|b1_q1|b1_q2|b1_q3|b1_q4|b1_q5|b1_q6|b1_q7 b1_c4_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3345 \$3043 a4|b0_p4|b1_p4|b2_p4|b3_p4|b4_p4|b5_p4|b6_p4|b7_p4 \$3324 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3346 b1_c4
+ b1_not|b1_q0_not|b1_q1_not|b1_q2_not|b1_q3_not|b1_q4_not|b1_q5_not|b1_q6_not|b1_q7_not
+ \$3043 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3347 \$3045
+ b0_not|b0_q0_not|b0_q1_not|b0_q3_not|b0_q4_not|b0_q5_not|b0_q6_not|b0_q7_not|b1_q2_not
+ b0_c5_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3348 \$3325 a5|b0_p5|b1_p5|b3_p5|b4_p5|b5_p5|b6_p5|b7_p5 \$3045 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3349 b0_c5 b0|b0_q0|b0_q1|b0_q2|b0_q3|b0_q4|b0_q5|b0_q6|b0_q7 \$3325 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3350 \$3327 b0|b0_q0|b0_q1|b0_q2|b0_q3|b0_q4|b0_q5|b0_q6|b0_q7 b0_c5_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3351 \$3047 a5|b0_p5|b1_p5|b3_p5|b4_p5|b5_p5|b6_p5|b7_p5 \$3327 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3352 b0_c5
+ b0_not|b0_q0_not|b0_q1_not|b0_q3_not|b0_q4_not|b0_q5_not|b0_q6_not|b0_q7_not|b1_q2_not
+ \$3047 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3353 \$3175 \$3047 \$3115 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3354 \$3177 \$3047 \$3043 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3355 \$3115 \$3045 \$3177 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3356 \$3176 \$3047 \$3116 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3357 \$3034 \$3047 \$3328 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3358 \$3116 \$3045 \$3034 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3359 \$3179 b0_r5_b \$3176 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3360 \$3181 \$3178 \$3175 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3361 \$3051
+ b2_not|b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not
+ b2_c4_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3362 \$3333 a4|b0_p4|b1_p4|b2_p4|b3_p4|b4_p4|b5_p4|b6_p4|b7_p4 \$3051 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3363 b2_c4 b2|b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7 \$3333 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3364 \$3334 b2|b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7 b2_c4_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3365 \$3053 a4|b0_p4|b1_p4|b2_p4|b3_p4|b4_p4|b5_p4|b6_p4|b7_p4 \$3334 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3366 b2_c4
+ b2_not|b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not
+ \$3053 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3367 \$3182 \$3053 \$2214 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3368 \$3184 \$3053 \$2213 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3369 \$2214 \$3051 \$3184 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3370 \$3183 \$3053 \$3117 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3371 \$3035 \$3053 \$3335 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3372 \$3117 \$3051 \$3035 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3373 \$3186 b2_r4_b \$3183 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3374 \$3188 \$3185 \$3182 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3375 \$3057
+ b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b3_not|b3_q0_not|b3_q1_not|b3_q2_not|b3_q3_not|b3_q4_not|b3_q5_not|b3_q6_not|b3_q7_not
+ b2_c4_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3376 \$3340 a4|b0_p4|b1_p4|b2_p4|b3_p4|b4_p4|b5_p4|b6_p4|b7_p4 \$3057 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3377 b2_c4
+ b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b3|b3_q0|b3_q1|b3_q2|b3_q3|b3_q4|b3_q5|b3_q6|b3_q7
+ \$3340 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3378 \$3341
+ b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b3|b3_q0|b3_q1|b3_q2|b3_q3|b3_q4|b3_q5|b3_q6|b3_q7
+ b2_c4_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3379 \$3058 a4|b0_p4|b1_p4|b2_p4|b3_p4|b4_p4|b5_p4|b6_p4|b7_p4 \$3341 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3380 b2_c4
+ b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b3_not|b3_q0_not|b3_q1_not|b3_q2_not|b3_q3_not|b3_q4_not|b3_q5_not|b3_q6_not|b3_q7_not
+ \$3058 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3381 \$2375 \$3191 \$3057 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3382 \$3343 \$3190 \$2375 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3383 \$3058 \$3189 \$3343 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3384 \$3344 \$3189 \$3057 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3385 \$2376 \$3190 \$3344 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3386 \$3058 \$3191 \$2376 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3387 b3_r4_b_not \$3191 \$2166 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3388 \$3345 \$3190 b3_r4_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3389 \$2165 \$3189 \$3345 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3390 \$3346 \$3189 \$2166 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3391 b3_r4_b \$3190 \$3346 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3392 \$2165 \$3191 b3_r4_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3393 \$3192 \$3064 \$2168 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3394 \$3194 \$3064 \$2167 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3395 \$3193 \$3064 \$3123 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3396 \$3037 \$3064 \$3349 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3397 b4_r4_b_not \$3194 \$2226 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3398 \$3352 \$3193 b4_r4_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3399 \$2225 \$3192 \$3352 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3400 \$3353 \$3192 \$2226 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3401 b4_r4_b \$3193 \$3353 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3402 \$2225 \$3194 b4_r4_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3403 \$3197 \$3070 \$2228 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3404 \$3199 \$3070 \$2227 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3405 \$3198 \$3070 \$3126 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3406 \$3038 \$3070 \$3356 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3407 b5_r4_b_not \$3199 \$2231 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3408 \$3359 \$3198 b5_r4_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3409 \$2230 \$3197 \$3359 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3410 \$3360 \$3197 \$2231 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3411 b5_r4_b \$3198 \$3360 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3412 \$2230 \$3199 b5_r4_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3413 \$3075
+ b6_not|b6_q0_not|b6_q1_not|b6_q2_not|b6_q3_not|b6_q4_not|b6_q5_not|b6_q6_not|b6_q7_not
+ b6_c4_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3414 \$3361 a4|b0_p4|b1_p4|b2_p4|b3_p4|b4_p4|b5_p4|b6_p4|b7_p4 \$3075 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3415 b6_c4 b6|b6_q0|b6_q1|b6_q2|b6_q3|b6_q4|b6_q5|b6_q6|b6_q7 \$3361 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3416 \$3363 b6|b6_q0|b6_q1|b6_q2|b6_q3|b6_q4|b6_q5|b6_q6|b6_q7 b6_c4_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3417 \$3077 a4|b0_p4|b1_p4|b2_p4|b3_p4|b4_p4|b5_p4|b6_p4|b7_p4 \$3363 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3418 b6_c4
+ b6_not|b6_q0_not|b6_q1_not|b6_q2_not|b6_q3_not|b6_q4_not|b6_q5_not|b6_q6_not|b6_q7_not
+ \$3077 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3419 \$3202 \$3077 \$2233 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3420 \$3204 \$3077 \$2232 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3421 \$3203 \$3077 \$3129 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3422 \$3039 \$3077 \$3364 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3423 b6_r4_b_not \$3204 \$2238 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3424 \$3367 \$3203 b6_r4_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3425 \$2237 \$3202 \$3367 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3426 \$3368 \$3202 \$2238 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3427 b6_r4_b \$3203 \$3368 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3428 \$2237 \$3204 b6_r4_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3429 \$3081
+ b7_not|b7_q0_not|b7_q1_not|b7_q2_not|b7_q3_not|b7_q4_not|b7_q5_not|b7_q6_not|b7_q7_not
+ \$3080 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3430 \$3369 a4|b0_p4|b1_p4|b2_p4|b3_p4|b4_p4|b5_p4|b6_p4|b7_p4 \$3081 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3431 \$3084 b1_q3|b7|b7_q0|b7_q1|b7_q2|b7_q4|b7_q5|b7_q6|b7_q7 \$3369 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3432 \$3370 b1_q3|b7|b7_q0|b7_q1|b7_q2|b7_q4|b7_q5|b7_q6|b7_q7 \$3080 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3433 \$3083 a4|b0_p4|b1_p4|b2_p4|b3_p4|b4_p4|b5_p4|b6_p4|b7_p4 \$3370 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3434 \$3084
+ b7_not|b7_q0_not|b7_q1_not|b7_q2_not|b7_q3_not|b7_q4_not|b7_q5_not|b7_q6_not|b7_q7_not
+ \$3083 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3435 \$3207 \$3083 \$2240 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3436 \$3209 \$3083 \$2239 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3437 \$3208 \$3083 \$3132 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3438 \$3040 \$3083 \$3371 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3439 \$3085 \$3209 \$2243 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3440 \$3374 \$3208 \$3085 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3441 \$2242 \$3207 \$3374 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3442 \$3375 \$3207 \$2243 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3443 \$3086 \$3208 \$3375 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3444 \$2242 \$3209 \$3086 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3445 \$4038
+ a3_not|b0_p3_not|b1_p3_not|b2_p3_not|b3_p3_not|b5_p3_not|b6_p3_not|b7_p3_not
+ b1_c3_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3446 b1_c3
+ a3_not|b0_p3_not|b1_p3_not|b2_p3_not|b3_p3_not|b5_p3_not|b6_p3_not|b7_p3_not
+ \$4039 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3447 \$4041
+ a4_not|b0_p4_not|b1_p4_not|b2_p4_not|b3_p4_not|b5_p4_not|b6_p4_not|b7_p4_not
+ b0_c4_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3448 b0_c4
+ a4_not|b0_p4_not|b1_p4_not|b2_p4_not|b3_p4_not|b5_p4_not|b6_p4_not|b7_p4_not
+ \$4042 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3449 \$2360 \$3177 \$3045 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3450 \$3329 \$3176 \$2360 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3451 \$3047 \$3175 \$3329 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3452 \$3330 \$3175 \$3045 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3453 \$2361 \$3176 \$3330 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3454 \$3047 \$3177 \$2361 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3455 b0_r5_b_not \$3177 \$2212 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3456 \$3331 \$3176 b0_r5_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3457 \$2211 \$3175 \$3331 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3458 \$3332 \$3175 \$2212 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3459 b0_r5_b \$3176 \$3332 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3460 \$2211 \$3177 b0_r5_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3461 \$2368 \$3184 \$3051 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3462 \$3336 \$3183 \$2368 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3463 \$3053 \$3182 \$3336 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3464 \$3337 \$3182 \$3051 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3465 \$2369 \$3183 \$3337 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3466 \$3053 \$3184 \$2369 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3467 b2_r4_b_not \$3184 \$2219 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3468 \$3338 \$3183 b2_r4_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3469 \$2218 \$3182 \$3338 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3470 \$3339 \$3182 \$2219 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3471 b2_r4_b \$3183 \$3339 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3472 \$2218 \$3184 b2_r4_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3473 \$4051
+ a3_not|b0_p3_not|b1_p3_not|b2_p3_not|b3_p3_not|b5_p3_not|b6_p3_not|b7_p3_not
+ b3_c2_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3474 b3_c2
+ a3_not|b0_p3_not|b1_p3_not|b2_p3_not|b3_p3_not|b5_p3_not|b6_p3_not|b7_p3_not
+ \$4052 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3475 \$3118 \$3620 \$4051 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3476 \$4052 \$3620 \$3342 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3477 b3_r3_b_not \$3620 \$3120 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3478 \$3119 \$3620 b3_r3_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3479 \$3062
+ b2_q0_not|b2_q1_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b4_not|b4_q7_not
+ b2_c4_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3480 \$3347 a4|b0_p4|b1_p4|b2_p4|b3_p4|b4_p4|b5_p4|b6_p4|b7_p4 \$3062 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3481 b2_c4 b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b4|b4_q7 \$3347 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3482 \$3348 b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b4|b4_q7 b2_c4_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3483 \$3064 a4|b0_p4|b1_p4|b2_p4|b3_p4|b4_p4|b5_p4|b6_p4|b7_p4 \$3348 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3484 b2_c4
+ b2_q0_not|b2_q1_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b4_not|b4_q7_not
+ \$3064 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3485 \$2383 \$3194 \$3062 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3486 \$3350 \$3193 \$2383 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3487 \$3064 \$3192 \$3350 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3488 \$3351 \$3192 \$3062 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3489 \$2384 \$3193 \$3351 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3490 \$3064 \$3194 \$2384 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3491 \$3068
+ b5_not|b5_q0_not|b5_q1_not|b5_q2_not|b5_q3_not|b5_q4_not|b5_q5_not|b5_q6_not|b5_q7_not
+ \$3067 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3492 \$3354 a4|b0_p4|b1_p4|b2_p4|b3_p4|b4_p4|b5_p4|b6_p4|b7_p4 \$3068 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3493 \$3071 b5|b5_q0|b5_q1|b5_q2|b5_q3|b5_q4|b5_q5|b5_q6|b5_q7 \$3354 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3494 \$3355 b5|b5_q0|b5_q1|b5_q2|b5_q3|b5_q4|b5_q5|b5_q6|b5_q7 \$3067 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3495 \$3070 a4|b0_p4|b1_p4|b2_p4|b3_p4|b4_p4|b5_p4|b6_p4|b7_p4 \$3355 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3496 \$3071
+ b5_not|b5_q0_not|b5_q1_not|b5_q2_not|b5_q3_not|b5_q4_not|b5_q5_not|b5_q6_not|b5_q7_not
+ \$3070 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3497 \$2391 \$3199 \$3068 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3498 \$3357 \$3198 \$2391 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3499 \$3070 \$3197 \$3357 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3500 \$3358 \$3197 \$3068 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3501 \$2392 \$3198 \$3358 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3502 \$3070 \$3199 \$2392 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3503 \$4066
+ a3_not|b0_p3_not|b1_p3_not|b2_p3_not|b3_p3_not|b5_p3_not|b6_p3_not|b7_p3_not
+ b6_c2_not|b6_c3_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3504 b6_c2|b6_c3
+ a3_not|b0_p3_not|b1_p3_not|b2_p3_not|b3_p3_not|b5_p3_not|b6_p3_not|b7_p3_not
+ \$4067 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3505 \$2398 \$3204 \$3075 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3506 \$3365 \$3203 \$2398 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3507 \$3077 \$3202 \$3365 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3508 \$3366 \$3202 \$3075 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3509 \$2399 \$3203 \$3366 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3510 \$3077 \$3204 \$2399 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3511 \$2406 \$3209 \$3081 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3512 \$3372 \$3208 \$2406 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3513 \$3083 \$3207 \$3372 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3514 \$3373 \$3207 \$3081 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3515 \$2407 \$3208 \$3373 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3516 \$3083 \$3209 \$2407 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3517 \$4046
+ a3_not|b0_p3_not|b1_p3_not|b2_p3_not|b3_p3_not|b5_p3_not|b6_p3_not|b7_p3_not
+ b2_c2_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3518 b2_c2
+ a3_not|b0_p3_not|b1_p3_not|b2_p3_not|b3_p3_not|b5_p3_not|b6_p3_not|b7_p3_not
+ \$4047 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3519 \$3123 \$3622 \$4056 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3520 \$4057 \$3622 \$3349 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3521 \$3126 \$3624 \$4061 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3522 \$4062 \$3624 \$3356 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3523 \$3129 \$3626 \$4066 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3524 \$4067 \$3626 \$3364 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3525 \$4071
+ a3_not|b0_p3_not|b1_p3_not|b2_p3_not|b3_p3_not|b5_p3_not|b6_p3_not|b7_p3_not
+ b6_c2_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3526 b6_c2
+ a3_not|b0_p3_not|b1_p3_not|b2_p3_not|b3_p3_not|b5_p3_not|b6_p3_not|b7_p3_not
+ \$4072 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3527 \$3132 \$3628 \$4071 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3528 \$4072 \$3628 \$3371 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3529 \$3116 \$3612 \$4041 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3530 \$4042 \$3612 \$3328 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3531 b0_r4_b_not \$3612 \$3179 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3532 \$3178 \$3612 b0_r4_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3533 \$3117 \$3616 \$4046 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3534 \$4047 \$3616 \$3335 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3535 b2_r3_b_not \$3616 \$3186 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3536 \$3185 \$3616 b2_r3_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3537 \$3187 \$4051 \$4087 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3538 \$3188 \$4051 \$4159 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3539 \$4309 \$4051 \$4088 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3540 \$4089 \$4051 \$3620 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3541 \$4056
+ a3_not|b0_p3_not|b1_p3_not|b2_p3_not|b3_p3_not|b5_p3_not|b6_p3_not|b7_p3_not
+ b4_c2_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3542 b4_c2
+ a3_not|b0_p3_not|b1_p3_not|b2_p3_not|b3_p3_not|b5_p3_not|b6_p3_not|b7_p3_not
+ \$4057 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3543 b4_r3_b_not \$3622 \$3124 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3544 \$3195 \$3622 b4_r3_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3545 \$4061
+ a3_not|b0_p3_not|b1_p3_not|b2_p3_not|b3_p3_not|b5_p3_not|b6_p3_not|b7_p3_not
+ b5_c2_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3546 b5_c2
+ a3_not|b0_p3_not|b1_p3_not|b2_p3_not|b3_p3_not|b5_p3_not|b6_p3_not|b7_p3_not
+ \$4062 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3547 b5_r3_b_not \$3624 \$3127 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3548 \$3200 \$3624 b5_r3_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3549 b6_r3_b_not \$3626 \$3130 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3550 \$3205 \$3626 b6_r3_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3551 \$4073 \$3628 \$3133 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3552 \$3210 \$3628 \$4074 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3553 \$4039 \$4041 \$4145 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3554 \$4038 \$4041 \$4147 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3555 \$4293 \$4041 \$4146 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3556 \$4085 \$4041 \$3612 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3557 \$3180 \$4046 \$4152 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3558 \$3181 \$4046 \$4154 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3559 \$4301 \$4046 \$4153 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3560 \$4086 \$4046 \$3616 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3561 \$4087 \$4052 \$3188 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3562 \$4159 \$4052 \$3187 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3563 \$4088 \$4052 \$4089 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3564 \$3620 \$4052 \$4309 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3565 \$4090 b3_r3_b \$3620 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3566 \$4088 b3_r3_b_not \$4090 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3567 \$4091 b3_r3_b \$4088 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3568 \$3620 b3_r3_b_not \$4091 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3569 \$4092 \$4090 \$4159 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3570 \$4087 \$4091 \$4092 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3571 \$4093 \$4090 \$4087 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3572 \$4159 \$4091 \$4093 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3573 \$4094 \$4057 \$3122 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3574 \$3121 \$4056 \$4094 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3575 \$3122 \$4056 \$4160 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3576 \$4095 \$4057 \$4096 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3577 \$4317 \$4056 \$4095 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3578 \$4096 \$4056 \$3622 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3579 \$4095 b4_r3_b_not \$4161 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3580 \$3622 b4_r3_b_not \$4162 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3581 \$4094 \$4162 \$4163 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3582 \$4160 \$4162 \$4164 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3583 \$4097 \$4062 \$3125 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3584 \$3196 \$4061 \$4097 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3585 \$3125 \$4061 \$4165 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3586 \$4098 \$4062 \$4099 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3587 \$4325 \$4061 \$4098 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3588 \$4099 \$4061 \$3624 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3589 \$4098 b5_r3_b_not \$4166 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3590 \$3624 b5_r3_b_not \$4167 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3591 \$4097 \$4167 \$4168 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3592 \$4165 \$4167 \$4169 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3593 \$4100 \$4067 \$3128 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3594 \$3201 \$4066 \$4100 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3595 \$3128 \$4066 \$4170 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3596 \$4101 \$4067 \$4102 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3597 \$4332 \$4066 \$4101 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3598 \$4102 \$4066 \$3626 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3599 \$4101 b6_r3_b_not \$4171 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3600 \$3626 b6_r3_b_not \$4172 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3601 \$4100 \$4172 \$4173 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3602 \$4170 \$4172 \$4174 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3603 \$4103 \$4072 \$3131 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3604 \$3206 \$4071 \$4103 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3605 \$3131 \$4071 \$4175 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3606 \$4104 \$4072 \$4105 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3607 \$4340 \$4071 \$4104 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3608 \$4105 \$4071 \$3628 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3609 \$4104 \$4073 \$4176 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3610 \$3628 \$4073 \$4177 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3611 \$4103 \$4177 p10 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3612 \$4175 \$4177 p10_not vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3613 \$4038
+ b1_not|b1_q0_not|b1_q1_not|b1_q2_not|b1_q3_not|b1_q4_not|b1_q5_not|b1_q6_not|b1_q7_not
+ b1_c3_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3614 \$4142 a3|b0_p3|b1_p3|b2_p3|b3_p3|b5_p3|b6_p3|b7_p3 \$4038 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3615 b1_c3 b1|b1_q0|b1_q1|b1_q2|b1_q3|b1_q4|b1_q5|b1_q6|b1_q7 \$4142 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3616 \$4144 b1|b1_q0|b1_q1|b1_q2|b1_q3|b1_q4|b1_q5|b1_q6|b1_q7 b1_c3_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3617 \$4039 a3|b0_p3|b1_p3|b2_p3|b3_p3|b5_p3|b6_p3|b7_p3 \$4144 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3618 b1_c3
+ b1_not|b1_q0_not|b1_q1_not|b1_q2_not|b1_q3_not|b1_q4_not|b1_q5_not|b1_q6_not|b1_q7_not
+ \$4039 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3619 \$4041
+ b0_not|b0_q0_not|b0_q1_not|b0_q3_not|b0_q4_not|b0_q5_not|b0_q6_not|b0_q7_not|b1_q2_not
+ b0_c4_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3620 \$4290 a4|b0_p4|b1_p4|b2_p4|b3_p4|b4_p4|b5_p4|b6_p4|b7_p4 \$4041 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3621 b0_c4 b0|b0_q0|b0_q1|b0_q2|b0_q3|b0_q4|b0_q5|b0_q6|b0_q7 \$4290 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3622 \$4292 b0|b0_q0|b0_q1|b0_q2|b0_q3|b0_q4|b0_q5|b0_q6|b0_q7 b0_c4_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3623 \$4042 a4|b0_p4|b1_p4|b2_p4|b3_p4|b4_p4|b5_p4|b6_p4|b7_p4 \$4292 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3624 b0_c4
+ b0_not|b0_q0_not|b0_q1_not|b0_q3_not|b0_q4_not|b0_q5_not|b0_q6_not|b0_q7_not|b1_q2_not
+ \$4042 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3625 \$4145 \$4042 \$4038 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3626 \$4147 \$4042 \$4039 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3627 \$4146 \$4042 \$4085 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3628 \$3612 \$4042 \$4293 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3629 \$4148 b0_r4_b \$3612 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3630 \$4146 b0_r4_b_not \$4148 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3631 \$4149 b0_r4_b \$4146 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3632 \$3612 b0_r4_b_not \$4149 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3633 \$4150 \$4148 \$4147 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3634 \$4145 \$4149 \$4150 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3635 \$4151 \$4148 \$4145 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3636 \$4147 \$4149 \$4151 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3637 \$4046
+ b2_not|b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not
+ b2_c2_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3638 \$4298 a3|b0_p3|b1_p3|b2_p3|b3_p3|b5_p3|b6_p3|b7_p3 \$4046 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3639 b2_c2 b2|b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7 \$4298 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3640 \$4300 b2|b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7 b2_c2_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3641 \$4047 a3|b0_p3|b1_p3|b2_p3|b3_p3|b5_p3|b6_p3|b7_p3 \$4300 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3642 b2_c2
+ b2_not|b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not
+ \$4047 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3643 \$4152 \$4047 \$3181 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3644 \$4154 \$4047 \$3180 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3645 \$4153 \$4047 \$4086 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3646 \$3616 \$4047 \$4301 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3647 \$4155 b2_r3_b \$3616 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3648 \$4153 b2_r3_b_not \$4155 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3649 \$4156 b2_r3_b \$4153 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3650 \$3616 b2_r3_b_not \$4156 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3651 \$4157 \$4155 \$4154 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3652 \$4152 \$4156 \$4157 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3653 \$4158 \$4155 \$4152 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3654 \$4154 \$4156 \$4158 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3655 \$4051
+ b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b3_not|b3_q0_not|b3_q1_not|b3_q2_not|b3_q3_not|b3_q4_not|b3_q5_not|b3_q6_not|b3_q7_not
+ b3_c2_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3656 \$4306 a3|b0_p3|b1_p3|b2_p3|b3_p3|b5_p3|b6_p3|b7_p3 \$4051 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3657 b3_c2
+ b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b3|b3_q0|b3_q1|b3_q2|b3_q3|b3_q4|b3_q5|b3_q6|b3_q7
+ \$4306 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3658 \$4308
+ b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b3|b3_q0|b3_q1|b3_q2|b3_q3|b3_q4|b3_q5|b3_q6|b3_q7
+ b3_c2_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3659 \$4052 a3|b0_p3|b1_p3|b2_p3|b3_p3|b5_p3|b6_p3|b7_p3 \$4308 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3660 b3_c2
+ b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b3_not|b3_q0_not|b3_q1_not|b3_q2_not|b3_q3_not|b3_q4_not|b3_q5_not|b3_q6_not|b3_q7_not
+ \$4052 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3661 \$3118 \$4159 \$4051 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3662 \$4310 \$4088 \$3118 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3663 \$4052 \$4087 \$4310 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3664 \$4311 \$4087 \$4051 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3665 \$3342 \$4088 \$4311 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3666 \$4052 \$4159 \$3342 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3667 b3_r3_b_not \$4159 \$3120 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3668 \$4312 \$4088 b3_r3_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3669 \$3119 \$4087 \$4312 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3670 \$4313 \$4087 \$3120 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3671 b3_r3_b \$4088 \$4313 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3672 \$3119 \$4159 b3_r3_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3673 \$4160 \$4057 \$3121 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3674 \$3622 \$4057 \$4317 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3675 \$3123 \$4160 \$4056 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3676 \$4318 \$4095 \$3123 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3677 \$4057 \$4094 \$4318 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3678 \$4319 \$4094 \$4056 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3679 \$3349 \$4095 \$4319 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3680 \$4057 \$4160 \$3349 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3681 \$4161 b4_r3_b \$3622 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3682 \$4162 b4_r3_b \$4095 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3683 \$4163 \$4161 \$4160 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3684 \$4164 \$4161 \$4094 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3685 \$4165 \$4062 \$3196 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3686 \$3624 \$4062 \$4325 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3687 \$3126 \$4165 \$4061 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3688 \$4326 \$4098 \$3126 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3689 \$4062 \$4097 \$4326 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3690 \$4327 \$4097 \$4061 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3691 \$3356 \$4098 \$4327 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3692 \$4062 \$4165 \$3356 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3693 \$4166 b5_r3_b \$3624 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3694 \$4167 b5_r3_b \$4098 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3695 \$4168 \$4166 \$4165 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3696 \$4169 \$4166 \$4097 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3697 \$4066
+ b6_not|b6_q0_not|b6_q1_not|b6_q2_not|b6_q3_not|b6_q4_not|b6_q5_not|b6_q6_not|b6_q7_not
+ b6_c2_not|b6_c3_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3698 \$4330 a3|b0_p3|b1_p3|b2_p3|b3_p3|b5_p3|b6_p3|b7_p3 \$4066 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3699 b6_c2|b6_c3 b6|b6_q0|b6_q1|b6_q2|b6_q3|b6_q4|b6_q5|b6_q6|b6_q7 \$4330
+ vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3700 \$4331 b6|b6_q0|b6_q1|b6_q2|b6_q3|b6_q4|b6_q5|b6_q6|b6_q7
+ b6_c2_not|b6_c3_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3701 \$4067 a3|b0_p3|b1_p3|b2_p3|b3_p3|b5_p3|b6_p3|b7_p3 \$4331 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3702 b6_c2|b6_c3
+ b6_not|b6_q0_not|b6_q1_not|b6_q2_not|b6_q3_not|b6_q4_not|b6_q5_not|b6_q6_not|b6_q7_not
+ \$4067 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3703 \$4170 \$4067 \$3201 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3704 \$3626 \$4067 \$4332 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3705 \$3129 \$4170 \$4066 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3706 \$4333 \$4101 \$3129 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3707 \$4067 \$4100 \$4333 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3708 \$4334 \$4100 \$4066 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3709 \$3364 \$4101 \$4334 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3710 \$4067 \$4170 \$3364 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3711 \$4171 b6_r3_b \$3626 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3712 \$4172 b6_r3_b \$4101 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3713 \$4173 \$4171 \$4170 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3714 \$4174 \$4171 \$4100 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3715 \$4071
+ b7_not|b7_q0_not|b7_q1_not|b7_q2_not|b7_q3_not|b7_q4_not|b7_q5_not|b7_q6_not|b7_q7_not
+ b6_c2_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3716 \$4337 a3|b0_p3|b1_p3|b2_p3|b3_p3|b5_p3|b6_p3|b7_p3 \$4071 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3717 b6_c2 b1_q3|b7|b7_q0|b7_q1|b7_q2|b7_q4|b7_q5|b7_q6|b7_q7 \$4337 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3718 \$4339 b1_q3|b7|b7_q0|b7_q1|b7_q2|b7_q4|b7_q5|b7_q6|b7_q7 b6_c2_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3719 \$4072 a3|b0_p3|b1_p3|b2_p3|b3_p3|b5_p3|b6_p3|b7_p3 \$4339 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3720 b6_c2
+ b7_not|b7_q0_not|b7_q1_not|b7_q2_not|b7_q3_not|b7_q4_not|b7_q5_not|b7_q6_not|b7_q7_not
+ \$4072 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3721 \$4175 \$4072 \$3206 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3722 \$3628 \$4072 \$4340 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3723 \$3132 \$4175 \$4071 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3724 \$4341 \$4104 \$3132 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3725 \$4072 \$4103 \$4341 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3726 \$4342 \$4103 \$4071 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3727 \$3371 \$4104 \$4342 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3728 \$4072 \$4175 \$3371 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3729 \$4176 \$4074 \$3628 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3730 \$4177 \$4074 \$4104 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3731 p10 \$4176 \$4175 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$3732 p10_not \$4176 \$4103 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3733 \$5255
+ a2_not|b0_p2_not|b1_p2_not|b2_p2_not|b3_p2_not|b5_p2_not|b6_p2_not|b7_p2_not
+ b1_c2_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3734 b1_c2
+ a2_not|b0_p2_not|b1_p2_not|b2_p2_not|b3_p2_not|b5_p2_not|b6_p2_not|b7_p2_not
+ \$5008 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3735 \$5010
+ a3_not|b0_p3_not|b1_p3_not|b2_p3_not|b3_p3_not|b5_p3_not|b6_p3_not|b7_p3_not
+ b0_c3_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3736 b0_c3
+ a3_not|b0_p3_not|b1_p3_not|b2_p3_not|b3_p3_not|b5_p3_not|b6_p3_not|b7_p3_not
+ \$5011 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3737 \$3116 \$4147 \$4041 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3738 \$4294 \$4146 \$3116 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3739 \$4042 \$4145 \$4294 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3740 \$4295 \$4145 \$4041 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3741 \$3328 \$4146 \$4295 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3742 \$4042 \$4147 \$3328 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3743 b0_r4_b_not \$4147 \$3179 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3744 \$4296 \$4146 b0_r4_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3745 \$3178 \$4145 \$4296 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3746 \$4297 \$4145 \$3179 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3747 b0_r4_b \$4146 \$4297 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3748 \$3178 \$4147 b0_r4_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3749 \$5015
+ a2_not|b0_p2_not|b1_p2_not|b2_p2_not|b3_p2_not|b5_p2_not|b6_p2_not|b7_p2_not
+ b2_c2_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3750 b2_c2
+ a2_not|b0_p2_not|b1_p2_not|b2_p2_not|b3_p2_not|b5_p2_not|b6_p2_not|b7_p2_not
+ \$5016 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3751 \$3117 \$4154 \$4046 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3752 \$4302 \$4153 \$3117 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3753 \$4047 \$4152 \$4302 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3754 \$4303 \$4152 \$4046 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3755 \$3335 \$4153 \$4303 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3756 \$4047 \$4154 \$3335 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3757 b2_r3_b_not \$4154 \$3186 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3758 \$4304 \$4153 b2_r3_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3759 \$3185 \$4152 \$4304 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3760 \$4305 \$4152 \$3186 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3761 b2_r3_b \$4153 \$4305 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3762 \$3185 \$4154 b2_r3_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3763 \$5020
+ a2_not|b0_p2_not|b1_p2_not|b2_p2_not|b3_p2_not|b5_p2_not|b6_p2_not|b7_p2_not
+ b3_c2_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3764 b3_c2
+ a2_not|b0_p2_not|b1_p2_not|b2_p2_not|b3_p2_not|b5_p2_not|b6_p2_not|b7_p2_not
+ \$5021 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3765 \$4056
+ b2_q0_not|b2_q1_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b4_not|b4_q7_not
+ b4_c2_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3766 \$4314 a3|b0_p3|b1_p3|b2_p3|b3_p3|b5_p3|b6_p3|b7_p3 \$4056 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3767 b4_c2 b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b4|b4_q7 \$4314 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3768 \$4316 b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b4|b4_q7 b4_c2_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3769 \$4057 a3|b0_p3|b1_p3|b2_p3|b3_p3|b5_p3|b6_p3|b7_p3 \$4316 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3770 b4_c2
+ b2_q0_not|b2_q1_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b4_not|b4_q7_not
+ \$4057 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3771 b4_r3_b_not \$4160 \$3124 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3772 \$4320 \$4095 b4_r3_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3773 \$3195 \$4094 \$4320 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3774 \$4321 \$4094 \$3124 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3775 b4_r3_b \$4095 \$4321 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3776 \$3195 \$4160 b4_r3_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3777 \$4061
+ b5_not|b5_q0_not|b5_q1_not|b5_q2_not|b5_q3_not|b5_q4_not|b5_q5_not|b5_q6_not|b5_q7_not
+ b5_c2_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3778 \$4322 a3|b0_p3|b1_p3|b2_p3|b3_p3|b5_p3|b6_p3|b7_p3 \$4061 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3779 b5_c2 b5|b5_q0|b5_q1|b5_q2|b5_q3|b5_q4|b5_q5|b5_q6|b5_q7 \$4322 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3780 \$4324 b5|b5_q0|b5_q1|b5_q2|b5_q3|b5_q4|b5_q5|b5_q6|b5_q7 b5_c2_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3781 \$4062 a3|b0_p3|b1_p3|b2_p3|b3_p3|b5_p3|b6_p3|b7_p3 \$4324 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3782 b5_c2
+ b5_not|b5_q0_not|b5_q1_not|b5_q2_not|b5_q3_not|b5_q4_not|b5_q5_not|b5_q6_not|b5_q7_not
+ \$4062 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3783 b5_r3_b_not \$4165 \$3127 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3784 \$4328 \$4098 b5_r3_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3785 \$3200 \$4097 \$4328 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3786 \$4329 \$4097 \$3127 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3787 b5_r3_b \$4098 \$4329 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3788 \$3200 \$4165 b5_r3_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3789 \$5035
+ a2_not|b0_p2_not|b1_p2_not|b2_p2_not|b3_p2_not|b5_p2_not|b6_p2_not|b7_p2_not
+ b6_c2_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3790 b6_c2
+ a2_not|b0_p2_not|b1_p2_not|b2_p2_not|b3_p2_not|b5_p2_not|b6_p2_not|b7_p2_not
+ \$5036 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3791 b6_r3_b_not \$4170 \$3130 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3792 \$4335 \$4101 b6_r3_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3793 \$3205 \$4100 \$4335 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3794 \$4336 \$4100 \$3130 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3795 b6_r3_b \$4101 \$4336 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3796 \$3205 \$4170 b6_r3_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3797 \$5040
+ a2_not|b0_p2_not|b1_p2_not|b2_p2_not|b3_p2_not|b5_p2_not|b6_p2_not|b7_p2_not
+ b6_c2_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3798 b6_c2
+ a2_not|b0_p2_not|b1_p2_not|b2_p2_not|b3_p2_not|b5_p2_not|b6_p2_not|b7_p2_not
+ \$5041 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3799 \$4073 \$4175 \$3133 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3800 \$4343 \$4104 \$4073 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3801 \$3210 \$4103 \$4343 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3802 \$4344 \$4103 \$3133 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3803 \$4074 \$4104 \$4344 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3804 \$3210 \$4175 \$4074 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3805 \$4089 \$4831 \$5020 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3806 \$5021 \$4831 \$4309 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3807 b3_r2_b_not \$4831 \$4091 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3808 \$4090 \$4831 b3_r2_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3809 \$5025
+ a2_not|b0_p2_not|b1_p2_not|b2_p2_not|b3_p2_not|b5_p2_not|b6_p2_not|b7_p2_not
+ b4_c2_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3810 b4_c2
+ a2_not|b0_p2_not|b1_p2_not|b2_p2_not|b3_p2_not|b5_p2_not|b6_p2_not|b7_p2_not
+ \$5026 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3811 b4_r2_b_not \$4835 \$4162 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3812 \$4161 \$4835 b4_r2_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3813 \$5030
+ a2_not|b0_p2_not|b1_p2_not|b2_p2_not|b3_p2_not|b5_p2_not|b6_p2_not|b7_p2_not
+ b5_c2_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3814 b5_c2
+ a2_not|b0_p2_not|b1_p2_not|b2_p2_not|b3_p2_not|b5_p2_not|b6_p2_not|b7_p2_not
+ \$5031 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3815 b5_r2_b_not \$4837 \$4167 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3816 \$4166 \$4837 b5_r2_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3817 b6_r2_b_not \$4839 \$4172 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3818 \$4171 \$4839 b6_r2_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3819 \$5042 \$4841 \$4177 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3820 \$4176 \$4841 \$5043 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3821 \$4085 \$4827 \$5010 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3822 \$5011 \$4827 \$4293 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3823 \$5012 \$4827 \$4149 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3824 \$4148 \$4827 \$5013 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3825 \$4086 \$4829 \$5015 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3826 \$5016 \$4829 \$4301 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3827 b2_r2_b_not \$4829 \$4156 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3828 \$4155 \$4829 b2_r2_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3829 \$4157 \$5020 \$5080 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3830 \$4158 \$5020 \$5081 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3831 \$5279 \$5020 \$5082 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3832 \$5278 \$5020 \$4831 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3833 \$5083 b3_r2_b \$4831 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3834 \$5082 b3_r2_b_not \$5083 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3835 \$5084 b3_r2_b \$5082 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3836 \$4831 b3_r2_b_not \$5084 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3837 \$5085 \$5083 \$5081 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3838 \$5080 \$5084 \$5085 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3839 \$5086 \$5083 \$5080 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3840 \$5081 \$5084 \$5086 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3841 \$4096 \$4835 \$5025 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3842 \$5026 \$4835 \$4317 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3843 \$4099 \$4837 \$5030 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3844 \$5031 \$4837 \$4325 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3845 \$4102 \$4839 \$5035 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3846 \$5036 \$4839 \$4332 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3847 \$4105 \$4841 \$5040 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3848 \$5041 \$4841 \$4340 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3849 \$5128 \$5012 \$5072 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3850 \$4827 \$5012 \$5073 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3851 \$5127 \$5073 \$5074 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3852 \$5261 \$5073 \$5075 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3853 \$5130 b2_r2_b_not \$5076 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3854 \$4829 b2_r2_b_not \$5077 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3855 \$5129 \$5077 \$5078 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3856 \$5272 \$5077 \$5079 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3857 \$5080 \$5021 \$4158 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3858 \$5081 \$5021 \$4157 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3859 \$5082 \$5021 \$5278 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3860 \$4831 \$5021 \$5279 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3861 \$4092 \$5025 \$5134 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3862 \$5290 \$5025 \$5135 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3863 \$5088 b4_r2_b \$4835 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3864 \$5135 b4_r2_b_not \$5088 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3865 \$4835 b4_r2_b_not \$5089 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3866 \$5090 \$5088 \$5087 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3867 \$5134 \$5089 \$5090 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3868 \$5087 \$5089 \$5091 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3869 \$4163 \$5030 \$5136 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3870 \$5300 \$5030 \$5137 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3871 \$5093 b5_r2_b \$4837 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3872 \$5137 b5_r2_b_not \$5093 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3873 \$4837 b5_r2_b_not \$5094 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3874 \$5095 \$5093 \$5092 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3875 \$5136 \$5094 \$5095 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3876 \$5092 \$5094 \$5096 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3877 \$4168 \$5035 \$5138 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3878 \$5309 \$5035 \$5139 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3879 \$5098 b6_r2_b \$4839 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3880 \$5139 b6_r2_b_not \$5098 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3881 \$4839 b6_r2_b_not \$5099 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3882 \$5100 \$5098 \$5097 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3883 \$5138 \$5099 \$5100 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3884 \$5097 \$5099 \$5101 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3885 \$4173 \$5040 \$5140 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3886 \$5319 \$5040 \$5141 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3887 \$5103 \$5043 \$4841 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3888 \$5141 \$5042 \$5103 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3889 \$4841 \$5042 \$5104 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3890 p9 \$5103 \$5102 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$3891 \$5140 \$5104 p9 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3892 \$5102 \$5104 p9_not vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3893 \$5255
+ b1_not|b1_q0_not|b1_q1_not|b1_q2_not|b1_q3_not|b1_q4_not|b1_q5_not|b1_q6_not|b1_q7_not
+ b1_c2_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3894 \$5123 a2|b0_p2|b1_p2|b2_p2|b3_p2|b4_p2|b5_p2|b6_p2|b7_p2 \$5255 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3895 b1_c2 b1|b1_q0|b1_q1|b1_q2|b1_q3|b1_q4|b1_q5|b1_q6|b1_q7 \$5123 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3896 \$5125 b1|b1_q0|b1_q1|b1_q2|b1_q3|b1_q4|b1_q5|b1_q6|b1_q7 b1_c2_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3897 \$5008 a2|b0_p2|b1_p2|b2_p2|b3_p2|b4_p2|b5_p2|b6_p2|b7_p2 \$5125 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3898 b1_c2
+ b1_not|b1_q0_not|b1_q1_not|b1_q2_not|b1_q3_not|b1_q4_not|b1_q5_not|b1_q6_not|b1_q7_not
+ \$5008 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3899 \$5010
+ b0_not|b0_q0_not|b0_q1_not|b0_q3_not|b0_q4_not|b0_q5_not|b0_q6_not|b0_q7_not|b1_q2_not
+ b0_c3_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3900 \$5257 a3|b0_p3|b1_p3|b2_p3|b3_p3|b5_p3|b6_p3|b7_p3 \$5010 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3901 b0_c3 b0|b0_q0|b0_q1|b0_q2|b0_q3|b0_q4|b0_q5|b0_q6|b0_q7 \$5257 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3902 \$5258 b0|b0_q0|b0_q1|b0_q2|b0_q3|b0_q4|b0_q5|b0_q6|b0_q7 b0_c3_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3903 \$5011 a3|b0_p3|b1_p3|b2_p3|b3_p3|b5_p3|b6_p3|b7_p3 \$5258 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3904 b0_c3
+ b0_not|b0_q0_not|b0_q1_not|b0_q3_not|b0_q4_not|b0_q5_not|b0_q6_not|b0_q7_not|b1_q2_not
+ \$5011 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3905 \$5127 \$5011 \$5255 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3906 \$5008 \$5010 \$5127 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3907 \$5261 \$5011 \$5008 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3908 \$5255 \$5010 \$5261 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3909 \$5128 \$5011 \$5259 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3910 \$5260 \$5010 \$5128 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3911 \$4827 \$5011 \$5260 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3912 \$5259 \$5010 \$4827 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3913 \$5072 \$5013 \$4827 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3914 \$5073 \$5013 \$5128 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3915 \$5074 \$5072 \$5261 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3916 \$5075 \$5072 \$5127 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3917 \$5129 \$5016 \$4151 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3918 \$4150 \$5015 \$5129 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3919 \$5272 \$5016 \$4150 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3920 \$4151 \$5015 \$5272 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3921 \$5130 \$5016 \$5270 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3922 \$5271 \$5015 \$5130 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$3923 \$4829 \$5016 \$5271 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3924 \$5270 \$5015 \$4829 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3925 \$5076 b2_r2_b \$4829 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3926 \$5077 b2_r2_b \$5130 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3927 \$5078 \$5076 \$5272 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3928 \$5079 \$5076 \$5129 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3929 \$5020
+ b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b3_not|b3_q0_not|b3_q1_not|b3_q2_not|b3_q3_not|b3_q4_not|b3_q5_not|b3_q6_not|b3_q7_not
+ b3_c2_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3930 \$5131 a2|b0_p2|b1_p2|b2_p2|b3_p2|b4_p2|b5_p2|b6_p2|b7_p2 \$5020 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3931 b3_c2
+ b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b3|b3_q0|b3_q1|b3_q2|b3_q3|b3_q4|b3_q5|b3_q6|b3_q7
+ \$5131 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3932 \$5133
+ b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b3|b3_q0|b3_q1|b3_q2|b3_q3|b3_q4|b3_q5|b3_q6|b3_q7
+ b3_c2_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3933 \$5021 a2|b0_p2|b1_p2|b2_p2|b3_p2|b4_p2|b5_p2|b6_p2|b7_p2 \$5133 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3934 b3_c2
+ b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b3_not|b3_q0_not|b3_q1_not|b3_q2_not|b3_q3_not|b3_q4_not|b3_q5_not|b3_q6_not|b3_q7_not
+ \$5021 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3935 \$5134 \$5026 \$4093 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3936 \$5087 \$5026 \$4092 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3937 \$4093 \$5025 \$5087 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3938 \$5135 \$5026 \$5289 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3939 \$4835 \$5026 \$5290 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3940 \$5289 \$5025 \$4835 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3941 \$5089 b4_r2_b \$5135 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3942 \$5091 \$5088 \$5134 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3943 \$5136 \$5031 \$4164 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3944 \$5092 \$5031 \$4163 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3945 \$4164 \$5030 \$5092 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3946 \$5137 \$5031 \$5299 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3947 \$4837 \$5031 \$5300 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3948 \$5299 \$5030 \$4837 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3949 \$5094 b5_r2_b \$5137 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3950 \$5096 \$5093 \$5136 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3951 \$5035
+ b6_not|b6_q0_not|b6_q1_not|b6_q2_not|b6_q3_not|b6_q4_not|b6_q5_not|b6_q6_not|b6_q7_not
+ b6_c2_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3952 \$5306 a2|b0_p2|b1_p2|b2_p2|b3_p2|b4_p2|b5_p2|b6_p2|b7_p2 \$5035 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3953 b6_c2 b6|b6_q0|b6_q1|b6_q2|b6_q3|b6_q4|b6_q5|b6_q6|b6_q7 \$5306 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3954 \$5307 b6|b6_q0|b6_q1|b6_q2|b6_q3|b6_q4|b6_q5|b6_q6|b6_q7 b6_c2_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3955 \$5036 a2|b0_p2|b1_p2|b2_p2|b3_p2|b4_p2|b5_p2|b6_p2|b7_p2 \$5307 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3956 b6_c2
+ b6_not|b6_q0_not|b6_q1_not|b6_q2_not|b6_q3_not|b6_q4_not|b6_q5_not|b6_q6_not|b6_q7_not
+ \$5036 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3957 \$5138 \$5036 \$4169 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3958 \$5097 \$5036 \$4168 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3959 \$4169 \$5035 \$5097 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3960 \$5139 \$5036 \$5308 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3961 \$4839 \$5036 \$5309 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3962 \$5308 \$5035 \$4839 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3963 \$5099 b6_r2_b \$5139 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3964 \$5101 \$5098 \$5138 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3965 \$5140 \$5041 \$4174 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3966 \$5102 \$5041 \$4173 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3967 \$4174 \$5040 \$5102 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3968 \$5141 \$5041 \$5318 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$3969 \$4841 \$5041 \$5319 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3970 \$5318 \$5040 \$4841 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$3971 \$5104 \$5043 \$5141 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3972 p9_not \$5103 \$5140 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$3973 \$5015
+ b2_not|b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not
+ b2_c2_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3974 \$5267 a2|b0_p2|b1_p2|b2_p2|b3_p2|b4_p2|b5_p2|b6_p2|b7_p2 \$5015 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3975 b2_c2 b2|b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7 \$5267 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3976 \$5269 b2|b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7 b2_c2_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3977 \$5016 a2|b0_p2|b1_p2|b2_p2|b3_p2|b4_p2|b5_p2|b6_p2|b7_p2 \$5269 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3978 b2_c2
+ b2_not|b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not
+ \$5016 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3979 b3_r2_b_not \$5081 \$4091 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3980 \$5282 \$5082 b3_r2_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3981 \$4090 \$5080 \$5282 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3982 \$5283 \$5080 \$4091 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$3983 b3_r2_b \$5082 \$5283 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3984 \$4090 \$5081 b3_r2_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$3985 \$5025
+ b2_q0_not|b2_q1_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b4_not|b4_q7_not
+ b4_c2_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3986 \$5285 a2|b0_p2|b1_p2|b2_p2|b3_p2|b4_p2|b5_p2|b6_p2|b7_p2 \$5025 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3987 b4_c2 b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b4|b4_q7 \$5285 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3988 \$5287 b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b4|b4_q7 b4_c2_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3989 \$5026 a2|b0_p2|b1_p2|b2_p2|b3_p2|b4_p2|b5_p2|b6_p2|b7_p2 \$5287 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3990 b4_c2
+ b2_q0_not|b2_q1_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b4_not|b4_q7_not
+ \$5026 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3991 \$5030
+ b5_not|b5_q0_not|b5_q1_not|b5_q2_not|b5_q3_not|b5_q4_not|b5_q5_not|b5_q6_not|b5_q7_not
+ b5_c2_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3992 \$5296 a2|b0_p2|b1_p2|b2_p2|b3_p2|b4_p2|b5_p2|b6_p2|b7_p2 \$5030 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3993 b5_c2 b5|b5_q0|b5_q1|b5_q2|b5_q3|b5_q4|b5_q5|b5_q6|b5_q7 \$5296 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3994 \$5298 b5|b5_q0|b5_q1|b5_q2|b5_q3|b5_q4|b5_q5|b5_q6|b5_q7 b5_c2_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3995 \$5031 a2|b0_p2|b1_p2|b2_p2|b3_p2|b4_p2|b5_p2|b6_p2|b7_p2 \$5298 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3996 b5_c2
+ b5_not|b5_q0_not|b5_q1_not|b5_q2_not|b5_q3_not|b5_q4_not|b5_q5_not|b5_q6_not|b5_q7_not
+ \$5031 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3997 \$5040
+ b7_not|b7_q0_not|b7_q1_not|b7_q2_not|b7_q3_not|b7_q4_not|b7_q5_not|b7_q6_not|b7_q7_not
+ b6_c2_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$3998 \$5315 a2|b0_p2|b1_p2|b2_p2|b3_p2|b4_p2|b5_p2|b6_p2|b7_p2 \$5040 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$3999 b6_c2 b1_q3|b7|b7_q0|b7_q1|b7_q2|b7_q4|b7_q5|b7_q6|b7_q7 \$5315 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4000 \$5317 b1_q3|b7|b7_q0|b7_q1|b7_q2|b7_q4|b7_q5|b7_q6|b7_q7 b6_c2_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4001 \$5041 a2|b0_p2|b1_p2|b2_p2|b3_p2|b4_p2|b5_p2|b6_p2|b7_p2 \$5317 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4002 b6_c2
+ b7_not|b7_q0_not|b7_q1_not|b7_q2_not|b7_q3_not|b7_q4_not|b7_q5_not|b7_q6_not|b7_q7_not
+ \$5041 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4003 \$5012 \$5261 \$4149 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4004 \$5264 \$5128 \$5012 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4005 \$4148 \$5127 \$5264 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4006 \$5265 \$5127 \$4149 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4007 \$5013 \$5128 \$5265 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4008 \$4148 \$5261 \$5013 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4009 b2_r2_b_not \$5272 \$4156 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4010 \$5275 \$5130 b2_r2_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4011 \$4155 \$5129 \$5275 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4012 \$5276 \$5129 \$4156 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4013 b2_r2_b \$5130 \$5276 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4014 \$4155 \$5272 b2_r2_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4015 \$4089 \$5081 \$5020 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4016 \$5280 \$5082 \$4089 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4017 \$5021 \$5080 \$5280 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4018 \$5281 \$5080 \$5020 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4019 \$4309 \$5082 \$5281 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4020 \$5021 \$5081 \$4309 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4021 \$4096 \$5087 \$5025 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4022 \$5291 \$5135 \$4096 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4023 \$5026 \$5134 \$5291 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4024 \$5292 \$5134 \$5025 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4025 \$4317 \$5135 \$5292 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4026 \$5026 \$5087 \$4317 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4027 b4_r2_b_not \$5087 \$4162 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4028 \$5293 \$5135 b4_r2_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4029 \$4161 \$5134 \$5293 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4030 \$5294 \$5134 \$4162 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4031 b4_r2_b \$5135 \$5294 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4032 \$4161 \$5087 b4_r2_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4033 \$4099 \$5092 \$5030 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4034 \$5301 \$5137 \$4099 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4035 \$5031 \$5136 \$5301 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4036 \$5302 \$5136 \$5030 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4037 \$4325 \$5137 \$5302 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4038 \$5031 \$5092 \$4325 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4039 b5_r2_b_not \$5092 \$4167 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4040 \$5303 \$5137 b5_r2_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4041 \$4166 \$5136 \$5303 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4042 \$5304 \$5136 \$4167 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4043 b5_r2_b \$5137 \$5304 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4044 \$4166 \$5092 b5_r2_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4045 \$4102 \$5097 \$5035 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4046 \$5310 \$5139 \$4102 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4047 \$5036 \$5138 \$5310 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4048 \$5311 \$5138 \$5035 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4049 \$4332 \$5139 \$5311 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4050 \$5036 \$5097 \$4332 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4051 b6_r2_b_not \$5097 \$4172 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4052 \$5312 \$5139 b6_r2_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4053 \$4171 \$5138 \$5312 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4054 \$5313 \$5138 \$4172 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4055 b6_r2_b \$5139 \$5313 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4056 \$4171 \$5097 b6_r2_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4057 \$4105 \$5102 \$5040 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4058 \$5320 \$5141 \$4105 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4059 \$5041 \$5140 \$5320 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4060 \$5321 \$5140 \$5040 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4061 \$4340 \$5141 \$5321 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4062 \$5041 \$5102 \$4340 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4063 \$5042 \$5102 \$4177 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4064 \$5322 \$5141 \$5042 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4065 \$4176 \$5140 \$5322 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4066 \$5323 \$5140 \$4177 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4067 \$5043 \$5141 \$5323 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4068 \$4176 \$5102 \$5043 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4069 \$6409
+ a1_not|b0_p1_not|b1_p1_not|b2_p1_not|b3_p1_not|b4_p1_not|b5_p1_not|b6_p1_not|b7_p1_not
+ b1_c1_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$4070 b1_c1
+ a1_not|b0_p1_not|b1_p1_not|b2_p1_not|b3_p1_not|b4_p1_not|b5_p1_not|b6_p1_not|b7_p1_not
+ \$5948 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4071 \$5995
+ a2_not|b0_p2_not|b1_p2_not|b2_p2_not|b3_p2_not|b5_p2_not|b6_p2_not|b7_p2_not
+ b0_c2_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$4072 b0_c2
+ a2_not|b0_p2_not|b1_p2_not|b2_p2_not|b3_p2_not|b5_p2_not|b6_p2_not|b7_p2_not
+ \$5996 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4073 \$5259 \$5798 \$5995 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4074 \$4085 \$5261 \$5010 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4075 \$5262 \$5128 \$4085 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4076 \$5011 \$5127 \$5262 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4077 \$5263 \$5127 \$5010 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4078 \$4293 \$5128 \$5263 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4079 \$5996 \$5798 \$5260 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4080 \$5011 \$5261 \$4293 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4081 \$5950 \$5798 \$5073 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4082 \$5072 \$5798 \$5951 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4083 \$6062 \$5951 \$5798 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4084 \$6061 \$5950 \$6062 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4085 \$6063 \$5951 \$6061 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4086 \$5798 \$5950 \$6063 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4087 \$6064 \$6062 \$6060 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4088 \$6059 \$6063 \$6064 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4089 \$6065 \$6062 \$6059 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4090 \$6060 \$6063 \$6065 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4091 \$5998
+ a1_not|b0_p1_not|b1_p1_not|b2_p1_not|b3_p1_not|b4_p1_not|b5_p1_not|b6_p1_not|b7_p1_not
+ b2_c1_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$4092 b2_c1
+ a1_not|b0_p1_not|b1_p1_not|b2_p1_not|b3_p1_not|b4_p1_not|b5_p1_not|b6_p1_not|b7_p1_not
+ \$5999 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4093 \$5270 \$5800 \$5998 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4094 \$4086 \$5272 \$5015 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4095 \$5273 \$5130 \$4086 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4096 \$5016 \$5129 \$5273 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4097 \$5274 \$5129 \$5015 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4098 \$4301 \$5130 \$5274 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4099 \$5999 \$5800 \$5271 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4100 \$5016 \$5272 \$4301 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4101 b2_r1_b_not \$5800 \$5077 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4102 \$5076 \$5800 b2_r1_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4103 \$6069 b2_r1_b \$5800 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4104 \$6068 b2_r1_b_not \$6069 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4105 \$6070 b2_r1_b \$6068 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4106 \$5800 b2_r1_b_not \$6070 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4107 \$6071 \$6069 \$6067 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4108 \$6066 \$6070 \$6071 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4109 \$6072 \$6069 \$6066 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4110 \$6067 \$6070 \$6072 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4111 \$5956
+ a1_not|b0_p1_not|b1_p1_not|b2_p1_not|b3_p1_not|b4_p1_not|b5_p1_not|b6_p1_not|b7_p1_not
+ b2_c1_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$4112 b3_c1
+ a1_not|b0_p1_not|b1_p1_not|b2_p1_not|b3_p1_not|b4_p1_not|b5_p1_not|b6_p1_not|b7_p1_not
+ \$6000 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4113 \$6073 \$6000 \$5079 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4114 \$5078 \$5956 \$6073 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4115 \$6074 \$6000 \$5078 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4116 \$5079 \$5956 \$6074 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4117 \$6075 \$6000 \$6180 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4118 \$6416 \$5956 \$6075 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4119 \$5802 \$6000 \$6416 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4120 \$6180 \$5956 \$5802 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4121 \$5278 \$5802 \$5956 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4122 \$6000 \$5802 \$5279 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4123 b3_r1_b_not \$5802 \$5084 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4124 \$5083 \$5802 b3_r1_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4125 \$6076 b3_r1_b \$5802 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4126 \$6075 b3_r1_b_not \$6076 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4127 \$6077 b3_r1_b \$6075 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4128 \$5802 b3_r1_b_not \$6077 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4129 \$6078 \$6076 \$6074 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4130 \$6073 \$6077 \$6078 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4131 \$6079 \$6076 \$6073 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4132 \$6074 \$6077 \$6079 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4133 \$6002
+ a1_not|b0_p1_not|b1_p1_not|b2_p1_not|b3_p1_not|b4_p1_not|b5_p1_not|b6_p1_not|b7_p1_not
+ b2_c1_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$4134 b4_c1
+ a1_not|b0_p1_not|b1_p1_not|b2_p1_not|b3_p1_not|b4_p1_not|b5_p1_not|b6_p1_not|b7_p1_not
+ \$6003 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4135 \$5289 \$5804 \$6002 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4136 \$6003 \$5804 \$5290 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4137 b4_r1_b_not \$5804 \$5089 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4138 \$5088 \$5804 b4_r1_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4139 \$6083 b4_r1_b \$5804 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4140 \$6082 b4_r1_b_not \$6083 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4141 \$6084 b4_r1_b \$6082 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4142 \$5804 b4_r1_b_not \$6084 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4143 \$6085 \$6083 \$6081 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4144 \$6080 \$6084 \$6085 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4145 \$6086 \$6083 \$6080 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4146 \$6081 \$6084 \$6086 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4147 \$6005
+ a1_not|b0_p1_not|b1_p1_not|b2_p1_not|b3_p1_not|b4_p1_not|b5_p1_not|b6_p1_not|b7_p1_not
+ \$6004 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4148 b5_c1
+ a1_not|b0_p1_not|b1_p1_not|b2_p1_not|b3_p1_not|b4_p1_not|b5_p1_not|b6_p1_not|b7_p1_not
+ \$6006 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4149 \$5299 \$5806 \$6005 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4150 \$6006 \$5806 \$5300 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4151 b5_r1_b_not \$5806 \$5094 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4152 \$5093 \$5806 b5_r1_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4153 \$6090 b5_r1_b \$5806 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4154 \$6089 b5_r1_b_not \$6090 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4155 \$6091 b5_r1_b \$6089 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4156 \$5806 b5_r1_b_not \$6091 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4157 \$6092 \$6090 \$6088 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4158 \$6087 \$6091 \$6092 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4159 \$6093 \$6090 \$6087 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4160 \$6088 \$6091 \$6093 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4161 \$6008
+ a1_not|b0_p1_not|b1_p1_not|b2_p1_not|b3_p1_not|b4_p1_not|b5_p1_not|b6_p1_not|b7_p1_not
+ b6_c1_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$4162 b6_c1
+ a1_not|b0_p1_not|b1_p1_not|b2_p1_not|b3_p1_not|b4_p1_not|b5_p1_not|b6_p1_not|b7_p1_not
+ \$6009 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4163 \$5308 \$5808 \$6008 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4164 \$6009 \$5808 \$5309 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4165 b6_r1_b_not \$5808 \$5099 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4166 \$5098 \$5808 b6_r1_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4167 \$6097 b6_r1_b \$5808 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4168 \$6096 b6_r1_b_not \$6097 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4169 \$6098 b6_r1_b \$6096 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4170 \$5808 b6_r1_b_not \$6098 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4171 \$6099 \$6097 \$6095 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4172 \$6094 \$6098 \$6099 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4173 \$6100 \$6097 \$6094 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4174 \$6095 \$6098 \$6100 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4175 \$6011
+ a1_not|b0_p1_not|b1_p1_not|b2_p1_not|b3_p1_not|b4_p1_not|b5_p1_not|b6_p1_not|b7_p1_not
+ \$6010 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4176 b6_c1
+ a1_not|b0_p1_not|b1_p1_not|b2_p1_not|b3_p1_not|b4_p1_not|b5_p1_not|b6_p1_not|b7_p1_not
+ \$6012 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4177 \$5318 \$5810 \$6011 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4178 \$6012 \$5810 \$5319 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4179 \$5970 \$5810 \$5104 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4180 \$5103 \$5810 \$5971 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4181 \$6104 \$5971 \$5810 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4182 \$6103 \$5970 \$6104 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4183 \$6105 \$5971 \$6103 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4184 \$5810 \$5970 \$6105 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4185 p8 \$6104 \$6102 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$4186 \$6101 \$6105 p8 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4187 p8_not \$6104 \$6101 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4188 \$6102 \$6105 p8_not vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4189 \$6409
+ b1_not|b1_q0_not|b1_q1_not|b1_q2_not|b1_q3_not|b1_q4_not|b1_q5_not|b1_q6_not|b1_q7_not
+ b1_c1_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$4190 \$6158 a1|b0_p1|b1_p1|b2_p1|b3_p1|b4_p1|b5_p1|b6_p1|b7_p1 \$6409 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4191 b1_c1 b1|b1_q0|b1_q1|b1_q2|b1_q3|b1_q4|b1_q5|b1_q6|b1_q7 \$6158 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4192 \$6160 b1|b1_q0|b1_q1|b1_q2|b1_q3|b1_q4|b1_q5|b1_q6|b1_q7 b1_c1_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4193 \$5948 a1|b0_p1|b1_p1|b2_p1|b3_p1|b4_p1|b5_p1|b6_p1|b7_p1 \$6160 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4194 b1_c1
+ b1_not|b1_q0_not|b1_q1_not|b1_q2_not|b1_q3_not|b1_q4_not|b1_q5_not|b1_q6_not|b1_q7_not
+ \$5948 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4195 \$6059 \$5996 \$6409 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4196 \$5948 \$5995 \$6059 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4197 \$6060 \$5996 \$5948 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4198 \$6409 \$5995 \$6060 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4199 \$6061 \$5996 \$6164 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4200 \$6411 \$5995 \$6061 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4201 \$5798 \$5996 \$6411 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4202 \$6164 \$5995 \$5798 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4203 \$5950 \$6060 \$5073 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4204 \$6167 \$6061 \$5950 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4205 \$5072 \$6059 \$6167 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4206 \$6168 \$6059 \$5073 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4207 \$5951 \$6061 \$6168 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4208 \$5072 \$6060 \$5951 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4209 \$6066 \$5999 \$5075 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4210 \$5074 \$5998 \$6066 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4211 \$6067 \$5999 \$5074 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4212 \$5075 \$5998 \$6067 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4213 \$6068 \$5999 \$6172 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4214 \$6413 \$5998 \$6068 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4215 \$5800 \$5999 \$6413 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4216 \$6172 \$5998 \$5800 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4217 b2_r1_b_not \$6067 \$5077 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4218 \$6175 \$6068 b2_r1_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4219 \$5076 \$6066 \$6175 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4220 \$6176 \$6066 \$5077 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4221 b2_r1_b \$6068 \$6176 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4222 \$5076 \$6067 b2_r1_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4223 b3_r1_b_not \$6074 \$5084 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4224 \$6183 \$6075 b3_r1_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4225 \$5083 \$6073 \$6183 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4226 \$6184 \$6073 \$5084 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4227 b3_r1_b \$6075 \$6184 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4228 \$5083 \$6074 b3_r1_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4229 \$6080 \$6003 \$5086 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4230 \$5085 \$6002 \$6080 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4231 \$6081 \$6003 \$5085 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4232 \$5086 \$6002 \$6081 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4233 \$6082 \$6003 \$6188 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4234 \$6419 \$6002 \$6082 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4235 \$5804 \$6003 \$6419 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4236 \$6188 \$6002 \$5804 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4237 b4_r1_b_not \$6081 \$5089 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4238 \$6191 \$6082 b4_r1_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4239 \$5088 \$6080 \$6191 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4240 \$6192 \$6080 \$5089 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4241 b4_r1_b \$6082 \$6192 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4242 \$5088 \$6081 b4_r1_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4243 \$6087 \$6006 \$5091 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4244 \$5090 \$6005 \$6087 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4245 \$6088 \$6006 \$5090 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4246 \$5091 \$6005 \$6088 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4247 \$6089 \$6006 \$6196 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4248 \$6422 \$6005 \$6089 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4249 \$5806 \$6006 \$6422 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4250 \$6196 \$6005 \$5806 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4251 b5_r1_b_not \$6088 \$5094 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4252 \$6199 \$6089 b5_r1_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4253 \$5093 \$6087 \$6199 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4254 \$6200 \$6087 \$5094 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4255 b5_r1_b \$6089 \$6200 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4256 \$5093 \$6088 b5_r1_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4257 \$6094 \$6009 \$5096 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4258 \$5095 \$6008 \$6094 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4259 \$6095 \$6009 \$5095 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4260 \$5096 \$6008 \$6095 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4261 \$6096 \$6009 \$6203 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4262 \$6425 \$6008 \$6096 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4263 \$5808 \$6009 \$6425 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4264 \$6203 \$6008 \$5808 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4265 b6_r1_b_not \$6095 \$5099 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4266 \$6206 \$6096 b6_r1_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4267 \$5098 \$6094 \$6206 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4268 \$6207 \$6094 \$5099 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4269 b6_r1_b \$6096 \$6207 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4270 \$5098 \$6095 b6_r1_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4271 \$6101 \$6012 \$5101 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4272 \$5100 \$6011 \$6101 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4273 \$6102 \$6012 \$5100 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4274 \$5101 \$6011 \$6102 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4275 \$6103 \$6012 \$6211 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4276 \$6427 \$6011 \$6103 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4277 \$5810 \$6012 \$6427 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4278 \$6211 \$6011 \$5810 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4279 \$5970 \$6102 \$5104 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4280 \$6214 \$6103 \$5970 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4281 \$5103 \$6101 \$6214 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4282 \$6215 \$6101 \$5104 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4283 \$5971 \$6103 \$6215 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4284 \$5103 \$6102 \$5971 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4285 \$5995
+ b0_not|b0_q0_not|b0_q1_not|b0_q3_not|b0_q4_not|b0_q5_not|b0_q6_not|b0_q7_not|b1_q2_not
+ b0_c2_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$4286 \$6161 a2|b0_p2|b1_p2|b2_p2|b3_p2|b4_p2|b5_p2|b6_p2|b7_p2 \$5995 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4287 b0_c2 b0|b0_q0|b0_q1|b0_q2|b0_q3|b0_q4|b0_q5|b0_q6|b0_q7 \$6161 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4288 \$6163 b0|b0_q0|b0_q1|b0_q2|b0_q3|b0_q4|b0_q5|b0_q6|b0_q7 b0_c2_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4289 \$5996 a2|b0_p2|b1_p2|b2_p2|b3_p2|b4_p2|b5_p2|b6_p2|b7_p2 \$6163 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4290 b0_c2
+ b0_not|b0_q0_not|b0_q1_not|b0_q3_not|b0_q4_not|b0_q5_not|b0_q6_not|b0_q7_not|b1_q2_not
+ \$5996 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4291 \$5259 \$6060 \$5995 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4292 \$6165 \$6061 \$5259 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4293 \$5996 \$6059 \$6165 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4294 \$6166 \$6059 \$5995 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4295 \$5260 \$6061 \$6166 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4296 \$5996 \$6060 \$5260 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4297 \$5270 \$6067 \$5998 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4298 \$6173 \$6068 \$5270 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4299 \$5999 \$6066 \$6173 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4300 \$6174 \$6066 \$5998 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4301 \$5271 \$6068 \$6174 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4302 \$5999 \$6067 \$5271 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4303 \$5956
+ b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b3_not|b3_q0_not|b3_q1_not|b3_q2_not|b3_q3_not|b3_q4_not|b3_q5_not|b3_q6_not|b3_q7_not
+ b2_c1_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$4304 \$6177 a1|b0_p1|b1_p1|b2_p1|b3_p1|b4_p1|b5_p1|b6_p1|b7_p1 \$5956 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4305 b3_c1
+ b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b3|b3_q0|b3_q1|b3_q2|b3_q3|b3_q4|b3_q5|b3_q6|b3_q7
+ \$6177 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4306 \$6179
+ b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b3|b3_q0|b3_q1|b3_q2|b3_q3|b3_q4|b3_q5|b3_q6|b3_q7
+ b2_c1_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$4307 \$6000 a1|b0_p1|b1_p1|b2_p1|b3_p1|b4_p1|b5_p1|b6_p1|b7_p1 \$6179 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4308 b3_c1
+ b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b3_not|b3_q0_not|b3_q1_not|b3_q2_not|b3_q3_not|b3_q4_not|b3_q5_not|b3_q6_not|b3_q7_not
+ \$6000 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4309 \$5278 \$6074 \$5956 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4310 \$6181 \$6075 \$5278 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4311 \$6000 \$6073 \$6181 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4312 \$6182 \$6073 \$5956 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4313 \$5279 \$6075 \$6182 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4314 \$6000 \$6074 \$5279 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4315 \$5289 \$6081 \$6002 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4316 \$6189 \$6082 \$5289 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4317 \$6003 \$6080 \$6189 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4318 \$6190 \$6080 \$6002 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4319 \$5290 \$6082 \$6190 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4320 \$6003 \$6081 \$5290 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4321 \$5299 \$6088 \$6005 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4322 \$6197 \$6089 \$5299 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4323 \$6006 \$6087 \$6197 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4324 \$6198 \$6087 \$6005 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4325 \$5300 \$6089 \$6198 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4326 \$6006 \$6088 \$5300 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4327 \$5308 \$6095 \$6008 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4328 \$6204 \$6096 \$5308 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4329 \$6009 \$6094 \$6204 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4330 \$6205 \$6094 \$6008 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4331 \$5309 \$6096 \$6205 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4332 \$6009 \$6095 \$5309 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4333 \$5318 \$6102 \$6011 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4334 \$6212 \$6103 \$5318 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4335 \$6012 \$6101 \$6212 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4336 \$6213 \$6101 \$6011 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4337 \$5319 \$6103 \$6213 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4338 \$6012 \$6102 \$5319 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4339 \$6929
+ a0_not|b0_p0_not|b1_p0_not|b2_p0_not|b3_p0_not|b5_p0_not|b6_p0_not|b7_p0_not
+ b1_c0_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$4340 b1_c0
+ a0_not|b0_p0_not|b1_p0_not|b2_p0_not|b3_p0_not|b5_p0_not|b6_p0_not|b7_p0_not
+ \$6930 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4341 \$7232
+ a1_not|b0_p1_not|b1_p1_not|b2_p1_not|b3_p1_not|b4_p1_not|b5_p1_not|b6_p1_not|b7_p1_not
+ b0_c1_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$4342 b0_c1
+ a1_not|b0_p1_not|b1_p1_not|b2_p1_not|b3_p1_not|b4_p1_not|b5_p1_not|b6_p1_not|b7_p1_not
+ \$6932 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4343 \$6164 \$6905 \$7232 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4344 \$6932 \$6905 \$6411 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4345 \$6933 \$6905 \$6063 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4346 \$6062 \$6905 \$6934 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4347 \$6999 \$6933 x0_c0_b vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4348 \$6997 x0_c0_b_not p1 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4349 \$5998
+ b2_not|b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not
+ b2_c1_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$4350 \$7238
+ a0_not|b0_p0_not|b1_p0_not|b2_p0_not|b3_p0_not|b5_p0_not|b6_p0_not|b7_p0_not
+ b2_c0_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$4351 \$6169 a1|b0_p1|b1_p1|b2_p1|b3_p1|b4_p1|b5_p1|b6_p1|b7_p1 \$5998 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4352 b2_c1 b2|b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7 \$6169 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4353 \$6171 b2|b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7 b2_c1_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4354 \$5999 a1|b0_p1|b1_p1|b2_p1|b3_p1|b4_p1|b5_p1|b6_p1|b7_p1 \$6171 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4355 b2_c1
+ b2_not|b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not
+ \$5999 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4356 b2_c0
+ a0_not|b0_p0_not|b1_p0_not|b2_p0_not|b3_p0_not|b5_p0_not|b6_p0_not|b7_p0_not
+ \$6936 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4357 \$6172 \$6907 \$7238 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4358 \$6936 \$6907 \$6413 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4359 b2_r0_b_not \$6907 \$6070 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4360 \$6069 \$6907 b2_r0_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4361 \$7006 b2_r0_b_not \$7007 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4362 \$7004 \$7008 p2 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4363 \$6940
+ a0_not|b0_p0_not|b1_p0_not|b2_p0_not|b3_p0_not|b5_p0_not|b6_p0_not|b7_p0_not
+ b2_c0_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$4364 b2_c0
+ a0_not|b0_p0_not|b1_p0_not|b2_p0_not|b3_p0_not|b5_p0_not|b6_p0_not|b7_p0_not
+ \$6941 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4365 \$6180 \$6908 \$6940 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4366 \$6941 \$6908 \$6416 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4367 b3_r0_b_not \$6908 \$6077 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4368 \$6076 \$6908 b3_r0_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4369 \$7014 b3_r0_b \$6908 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4370 \$7013 b3_r0_b_not \$7014 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4371 \$7015 b3_r0_b \$7013 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4372 \$6908 b3_r0_b_not \$7015 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4373 p3 \$7014 \$7012 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$4374 \$7011 \$7015 p3 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4375 p3_not \$7014 \$7011 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4376 \$7012 \$7015 p3_not vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4377 \$6002
+ b2_q0_not|b2_q1_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b4_not|b4_q7_not
+ b2_c1_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$4378 \$7248
+ a0_not|b0_p0_not|b1_p0_not|b2_p0_not|b3_p0_not|b5_p0_not|b6_p0_not|b7_p0_not
+ b2_c0_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$4379 \$6185 a1|b0_p1|b1_p1|b2_p1|b3_p1|b4_p1|b5_p1|b6_p1|b7_p1 \$6002 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4380 b4_c1 b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b4|b4_q7 \$6185 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4381 \$6187 b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b4|b4_q7 b2_c1_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4382 \$6003 a1|b0_p1|b1_p1|b2_p1|b3_p1|b4_p1|b5_p1|b6_p1|b7_p1 \$6187 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4383 b4_c1
+ b2_q0_not|b2_q1_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b4_not|b4_q7_not
+ \$6003 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4384 b2_c0
+ a0_not|b0_p0_not|b1_p0_not|b2_p0_not|b3_p0_not|b5_p0_not|b6_p0_not|b7_p0_not
+ \$6945 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4385 \$6188 \$6909 \$7248 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4386 \$6945 \$6909 \$6419 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4387 b4_r0_b_not \$6909 \$6084 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4388 \$6083 \$6909 b4_r0_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4389 \$7020 b4_r0_b_not \$7021 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4390 \$6909 b4_r0_b_not \$7022 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4391 \$7018 \$7022 p4 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4392 \$7019 \$7022 p4_not vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4393 \$6005
+ b5_not|b5_q0_not|b5_q1_not|b5_q2_not|b5_q3_not|b5_q4_not|b5_q5_not|b5_q6_not|b5_q7_not
+ \$6004 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4394 \$7254
+ a0_not|b0_p0_not|b1_p0_not|b2_p0_not|b3_p0_not|b5_p0_not|b6_p0_not|b7_p0_not
+ \$6948 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4395 \$6193 a1|b0_p1|b1_p1|b2_p1|b3_p1|b4_p1|b5_p1|b6_p1|b7_p1 \$6005 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4396 b5_c1 b5|b5_q0|b5_q1|b5_q2|b5_q3|b5_q4|b5_q5|b5_q6|b5_q7 \$6193 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4397 \$6195 b5|b5_q0|b5_q1|b5_q2|b5_q3|b5_q4|b5_q5|b5_q6|b5_q7 \$6004 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4398 \$6006 a1|b0_p1|b1_p1|b2_p1|b3_p1|b4_p1|b5_p1|b6_p1|b7_p1 \$6195 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4399 b5_c1
+ b5_not|b5_q0_not|b5_q1_not|b5_q2_not|b5_q3_not|b5_q4_not|b5_q5_not|b5_q6_not|b5_q7_not
+ \$6006 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4400 \$6950
+ a0_not|b0_p0_not|b1_p0_not|b2_p0_not|b3_p0_not|b5_p0_not|b6_p0_not|b7_p0_not
+ \$6949 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4401 \$6196 \$6910 \$7254 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4402 \$6949 \$6910 \$6422 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4403 b5_r0_b_not \$6910 \$6091 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4404 \$6090 \$6910 b5_r0_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4405 \$7027 b5_r0_b_not \$7028 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4406 \$6910 b5_r0_b_not \$7029 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4407 \$7025 \$7029 p5 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4408 \$7026 \$7029 p5_not vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4409 \$6008
+ b6_not|b6_q0_not|b6_q1_not|b6_q2_not|b6_q3_not|b6_q4_not|b6_q5_not|b6_q6_not|b6_q7_not
+ b6_c1_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$4410 \$7261
+ a0_not|b0_p0_not|b1_p0_not|b2_p0_not|b3_p0_not|b5_p0_not|b6_p0_not|b7_p0_not
+ b6_c0_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$4411 \$6201 a1|b0_p1|b1_p1|b2_p1|b3_p1|b4_p1|b5_p1|b6_p1|b7_p1 \$6008 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4412 b6_c1 b6|b6_q0|b6_q1|b6_q2|b6_q3|b6_q4|b6_q5|b6_q6|b6_q7 \$6201 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4413 \$6202 b6|b6_q0|b6_q1|b6_q2|b6_q3|b6_q4|b6_q5|b6_q6|b6_q7 b6_c1_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4414 \$6009 a1|b0_p1|b1_p1|b2_p1|b3_p1|b4_p1|b5_p1|b6_p1|b7_p1 \$6202 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4415 b6_c1
+ b6_not|b6_q0_not|b6_q1_not|b6_q2_not|b6_q3_not|b6_q4_not|b6_q5_not|b6_q6_not|b6_q7_not
+ \$6009 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4416 b6_c0
+ a0_not|b0_p0_not|b1_p0_not|b2_p0_not|b3_p0_not|b5_p0_not|b6_p0_not|b7_p0_not
+ \$6954 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4417 \$6203 \$6911 \$7261 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4418 \$6954 \$6911 \$6425 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4419 b6_r0_b_not \$6911 \$6098 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4420 \$6097 \$6911 b6_r0_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4421 \$7034 b6_r0_b_not \$7035 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4422 \$6911 b6_r0_b_not \$7036 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4423 \$7032 \$7036 p6 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4424 \$7033 \$7036 p6_not vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4425 \$6011
+ b7_not|b7_q0_not|b7_q1_not|b7_q2_not|b7_q3_not|b7_q4_not|b7_q5_not|b7_q6_not|b7_q7_not
+ \$6010 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4426 \$7267
+ a0_not|b0_p0_not|b1_p0_not|b2_p0_not|b3_p0_not|b5_p0_not|b6_p0_not|b7_p0_not
+ \$6957 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4427 \$6208 a1|b0_p1|b1_p1|b2_p1|b3_p1|b4_p1|b5_p1|b6_p1|b7_p1 \$6011 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4428 b6_c1 b1_q3|b7|b7_q0|b7_q1|b7_q2|b7_q4|b7_q5|b7_q6|b7_q7 \$6208 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4429 \$6210 b1_q3|b7|b7_q0|b7_q1|b7_q2|b7_q4|b7_q5|b7_q6|b7_q7 \$6010 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4430 \$6012 a1|b0_p1|b1_p1|b2_p1|b3_p1|b4_p1|b5_p1|b6_p1|b7_p1 \$6210 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4431 b6_c1
+ b7_not|b7_q0_not|b7_q1_not|b7_q2_not|b7_q3_not|b7_q4_not|b7_q5_not|b7_q6_not|b7_q7_not
+ \$6012 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4432 \$6959
+ a0_not|b0_p0_not|b1_p0_not|b2_p0_not|b3_p0_not|b5_p0_not|b6_p0_not|b7_p0_not
+ \$6958 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4433 \$6211 \$6912 \$7267 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4434 \$6958 \$6912 \$6427 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4435 \$6960 \$6912 \$6105 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4436 \$6104 \$6912 \$6961 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4437 \$7041 \$6960 \$7042 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4438 \$6912 \$6960 \$7043 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4439 \$7039 \$7043 p7 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4440 \$7040 \$7043 p7_not vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4441 \$6930 \$7232 \$6997 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4442 \$6929 \$7232 \$6998 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4443 x0_c0_f \$7232 \$6999 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4444 x0_c0_f_not \$7232 \$6905 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4445 x0_c0_b \$6934 \$6905 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4446 x0_c0_b_not \$6934 \$6999 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4447 \$6905 \$6933 x0_c0_b_not vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4448 p1 x0_c0_b \$6998 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$4449 p1_not x0_c0_b \$6997 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4450 \$6998 x0_c0_b_not p1_not vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4451 \$6064 \$7238 \$7004 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4452 \$6065 \$7238 \$7005 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4453 \$7080 \$7238 \$7006 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4454 \$7239 \$7238 \$6907 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4455 \$7007 b2_r0_b \$6907 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4456 \$7008 b2_r0_b \$7006 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4457 \$6907 b2_r0_b_not \$7008 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4458 p2 \$7007 \$7005 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$4459 p2_not \$7007 \$7004 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4460 \$7005 \$7008 p2_not vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4461 \$7011 \$6941 \$6072 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4462 \$6071 \$6940 \$7011 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4463 \$7012 \$6941 \$6071 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4464 \$6072 \$6940 \$7012 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4465 \$7013 \$6941 \$7242 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4466 \$7088 \$6940 \$7013 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4467 \$6908 \$6941 \$7088 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4468 \$7242 \$6940 \$6908 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4469 \$7018 \$6945 \$6079 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4470 \$6078 \$7248 \$7018 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4471 \$7019 \$6945 \$6078 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4472 \$6079 \$7248 \$7019 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4473 \$7020 \$6945 \$7249 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4474 \$7093 \$7248 \$7020 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4475 \$6909 \$6945 \$7093 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4476 \$7249 \$7248 \$6909 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4477 \$7021 b4_r0_b \$6909 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4478 \$7022 b4_r0_b \$7020 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4479 p4 \$7021 \$7019 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$4480 p4_not \$7021 \$7018 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4481 \$7025 \$6949 \$6086 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4482 \$6085 \$7254 \$7025 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4483 \$7026 \$6949 \$6085 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4484 \$6086 \$7254 \$7026 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4485 \$7027 \$6949 \$7255 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4486 \$7098 \$7254 \$7027 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4487 \$6910 \$6949 \$7098 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4488 \$7255 \$7254 \$6910 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4489 \$7028 b5_r0_b \$6910 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4490 \$7029 b5_r0_b \$7027 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4491 p5 \$7028 \$7026 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$4492 p5_not \$7028 \$7025 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4493 \$7032 \$6954 \$6093 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4494 \$6092 \$7261 \$7032 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4495 \$7033 \$6954 \$6092 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4496 \$6093 \$7261 \$7033 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4497 \$7034 \$6954 \$7262 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4498 \$7103 \$7261 \$7034 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4499 \$6911 \$6954 \$7103 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4500 \$7262 \$7261 \$6911 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4501 \$7035 b6_r0_b \$6911 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4502 \$7036 b6_r0_b \$7034 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4503 p6 \$7035 \$7033 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$4504 p6_not \$7035 \$7032 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4505 \$7039 \$6958 \$6100 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4506 \$6099 \$7267 \$7039 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4507 \$7040 \$6958 \$6099 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4508 \$6100 \$7267 \$7040 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4509 \$7041 \$6958 \$7268 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4510 \$7108 \$7267 \$7041 vss nfet_03v3 L=0.55U W=1.415U AS=0.742875P
+ AD=0.657975P PS=3.88U PD=3.76U
M$4511 \$6912 \$6958 \$7108 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4512 \$7268 \$7267 \$6912 vss nfet_03v3 L=0.55U W=1.385U AS=0.671725P
+ AD=0.6925P PS=3.74U PD=3.77U
M$4513 \$7042 \$6961 \$6912 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4514 \$7043 \$6961 \$7041 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4515 p7 \$7042 \$7040 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P AD=0.6576P
+ PS=3.67U PD=3.7U
M$4516 p7_not \$7042 \$7039 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4517 \$6929
+ b1_not|b1_q0_not|b1_q1_not|b1_q2_not|b1_q3_not|b1_q4_not|b1_q5_not|b1_q6_not|b1_q7_not
+ b1_c0_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$4518 \$7072 a0|b0_p0|b1_p0|b2_p0|b3_p0|b4_p0|b5_p0|b6_p0|b7_p0 \$6929 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4519 b1_c0 b1|b1_q0|b1_q1|b1_q2|b1_q3|b1_q4|b1_q5|b1_q6|b1_q7 \$7072 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4520 \$7074 b1|b1_q0|b1_q1|b1_q2|b1_q3|b1_q4|b1_q5|b1_q6|b1_q7 b1_c0_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4521 \$6930 a0|b0_p0|b1_p0|b2_p0|b3_p0|b4_p0|b5_p0|b6_p0|b7_p0 \$7074 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4522 b1_c0
+ b1_not|b1_q0_not|b1_q1_not|b1_q2_not|b1_q3_not|b1_q4_not|b1_q5_not|b1_q6_not|b1_q7_not
+ \$6930 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4523 \$7232
+ b0_not|b0_q0_not|b0_q1_not|b0_q3_not|b0_q4_not|b0_q5_not|b0_q6_not|b0_q7_not|b1_q2_not
+ b0_c1_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$4524 \$7227 a1|b0_p1|b1_p1|b2_p1|b3_p1|b4_p1|b5_p1|b6_p1|b7_p1 \$7232 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4525 b0_c1 b0|b0_q0|b0_q1|b0_q2|b0_q3|b0_q4|b0_q5|b0_q6|b0_q7 \$7227 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4526 \$7228 b0|b0_q0|b0_q1|b0_q2|b0_q3|b0_q4|b0_q5|b0_q6|b0_q7 b0_c1_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4527 \$6932 a1|b0_p1|b1_p1|b2_p1|b3_p1|b4_p1|b5_p1|b6_p1|b7_p1 \$7228 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4528 b0_c1
+ b0_not|b0_q0_not|b0_q1_not|b0_q3_not|b0_q4_not|b0_q5_not|b0_q6_not|b0_q7_not|b1_q2_not
+ \$6932 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4529 \$6997 \$6932 \$6929 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4530 \$6998 \$6932 \$6930 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4531 \$6999 \$6932 x0_c0_f_not vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4532 \$6905 \$6932 x0_c0_f vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4533 \$6164 \$6998 \$7232 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4534 \$7076 \$6999 \$6164 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4535 \$6932 \$6997 \$7076 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4536 \$7077 \$6997 \$7232 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4537 \$6411 \$6999 \$7077 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4538 \$6932 \$6998 \$6411 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4539 \$6933 \$6998 \$6063 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4540 \$7078 \$6999 \$6933 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4541 \$6062 \$6997 \$7078 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4542 \$7079 \$6997 \$6063 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4543 \$6934 \$6999 \$7079 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4544 \$6062 \$6998 \$6934 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4545 \$7238
+ b2_not|b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not
+ b2_c0_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$4546 \$7234 a0|b0_p0|b1_p0|b2_p0|b3_p0|b4_p0|b5_p0|b6_p0|b7_p0 \$7238 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4547 b2_c0 b2|b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7 \$7234 vss nfet_03v3
+ L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4548 \$7236 b2|b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7 b2_c0_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4549 \$6936 a0|b0_p0|b1_p0|b2_p0|b3_p0|b4_p0|b5_p0|b6_p0|b7_p0 \$7236 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4550 b2_c0
+ b2_not|b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not
+ \$6936 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4551 \$7004 \$6936 \$6065 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4552 \$7005 \$6936 \$6064 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4553 \$7006 \$6936 \$7239 vss nfet_03v3 L=0.55U W=1.37U AS=0.63705P
+ AD=0.6576P PS=3.67U PD=3.7U
M$4554 \$6907 \$6936 \$7080 vss nfet_03v3 L=0.55U W=1.365U AS=0.648375P
+ AD=0.64155P PS=3.68U PD=3.67U
M$4555 \$6172 \$7005 \$7238 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4556 \$7081 \$7006 \$6172 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4557 \$6936 \$7004 \$7081 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4558 \$7082 \$7004 \$7238 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4559 \$6413 \$7006 \$7082 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4560 \$6936 \$7005 \$6413 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4561 b2_r0_b_not \$7005 \$6070 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4562 \$7083 \$7006 b2_r0_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4563 \$6069 \$7004 \$7083 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4564 \$7084 \$7004 \$6070 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4565 b2_r0_b \$7006 \$7084 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4566 \$6069 \$7005 b2_r0_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4567 \$6940
+ b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b3_not|b3_q0_not|b3_q1_not|b3_q2_not|b3_q3_not|b3_q4_not|b3_q5_not|b3_q6_not|b3_q7_not
+ b2_c0_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$4568 \$7085 a0|b0_p0|b1_p0|b2_p0|b3_p0|b4_p0|b5_p0|b6_p0|b7_p0 \$6940 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4569 b2_c0
+ b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b3|b3_q0|b3_q1|b3_q2|b3_q3|b3_q4|b3_q5|b3_q6|b3_q7
+ \$7085 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4570 \$7087
+ b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b3|b3_q0|b3_q1|b3_q2|b3_q3|b3_q4|b3_q5|b3_q6|b3_q7
+ b2_c0_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$4571 \$6941 a0|b0_p0|b1_p0|b2_p0|b3_p0|b4_p0|b5_p0|b6_p0|b7_p0 \$7087 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4572 b2_c0
+ b2_q0_not|b2_q1_not|b2_q2_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b3_not|b3_q0_not|b3_q1_not|b3_q2_not|b3_q3_not|b3_q4_not|b3_q5_not|b3_q6_not|b3_q7_not
+ \$6941 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4573 \$6180 \$7012 \$6940 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4574 \$7089 \$7013 \$6180 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4575 \$6941 \$7011 \$7089 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4576 \$7090 \$7011 \$6940 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4577 \$6416 \$7013 \$7090 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4578 \$6941 \$7012 \$6416 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4579 b3_r0_b_not \$7012 \$6077 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4580 \$7091 \$7013 b3_r0_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4581 \$6076 \$7011 \$7091 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4582 \$7092 \$7011 \$6077 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4583 b3_r0_b \$7013 \$7092 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4584 \$6076 \$7012 b3_r0_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4585 \$7248
+ b2_q0_not|b2_q1_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b4_not|b4_q7_not
+ b2_c0_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$4586 \$7244 a0|b0_p0|b1_p0|b2_p0|b3_p0|b4_p0|b5_p0|b6_p0|b7_p0 \$7248 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4587 b2_c0 b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b4|b4_q7 \$7244 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4588 \$7246 b2_q0|b2_q1|b2_q2|b2_q3|b2_q4|b2_q5|b2_q7|b4|b4_q7 b2_c0_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4589 \$6945 a0|b0_p0|b1_p0|b2_p0|b3_p0|b4_p0|b5_p0|b6_p0|b7_p0 \$7246 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4590 b2_c0
+ b2_q0_not|b2_q1_not|b2_q3_not|b2_q4_not|b2_q5_not|b2_q7_not|b4_not|b4_q7_not
+ \$6945 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4591 \$6188 \$7019 \$7248 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4592 \$7094 \$7020 \$6188 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4593 \$6945 \$7018 \$7094 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4594 \$7095 \$7018 \$7248 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4595 \$6419 \$7020 \$7095 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4596 \$6945 \$7019 \$6419 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4597 b4_r0_b_not \$7019 \$6084 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4598 \$7096 \$7020 b4_r0_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4599 \$6083 \$7018 \$7096 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4600 \$7097 \$7018 \$6084 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4601 b4_r0_b \$7020 \$7097 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4602 \$6083 \$7019 b4_r0_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4603 \$6196 \$7026 \$7254 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4604 \$7099 \$7027 \$6196 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4605 \$6949 \$7025 \$7099 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4606 \$7100 \$7025 \$7254 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4607 \$6422 \$7027 \$7100 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4608 \$6949 \$7026 \$6422 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4609 b5_r0_b_not \$7026 \$6091 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4610 \$7101 \$7027 b5_r0_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4611 \$6090 \$7025 \$7101 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4612 \$7102 \$7025 \$6091 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4613 b5_r0_b \$7027 \$7102 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4614 \$6090 \$7026 b5_r0_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4615 \$7261
+ b6_not|b6_q0_not|b6_q1_not|b6_q2_not|b6_q3_not|b6_q4_not|b6_q5_not|b6_q6_not|b6_q7_not
+ b6_c0_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$4616 \$7257 a0|b0_p0|b1_p0|b2_p0|b3_p0|b4_p0|b5_p0|b6_p0|b7_p0 \$7261 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4617 b6_c0 b6|b6_q0|b6_q1|b6_q2|b6_q3|b6_q4|b6_q5|b6_q6|b6_q7 \$7257 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4618 \$7259 b6|b6_q0|b6_q1|b6_q2|b6_q3|b6_q4|b6_q5|b6_q6|b6_q7 b6_c0_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4619 \$6954 a0|b0_p0|b1_p0|b2_p0|b3_p0|b4_p0|b5_p0|b6_p0|b7_p0 \$7259 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4620 b6_c0
+ b6_not|b6_q0_not|b6_q1_not|b6_q2_not|b6_q3_not|b6_q4_not|b6_q5_not|b6_q6_not|b6_q7_not
+ \$6954 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4621 \$6203 \$7033 \$7261 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4622 \$7104 \$7034 \$6203 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4623 \$6954 \$7032 \$7104 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4624 \$7105 \$7032 \$7261 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4625 \$6425 \$7034 \$7105 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4626 \$6954 \$7033 \$6425 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4627 b6_r0_b_not \$7033 \$6098 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4628 \$7106 \$7034 b6_r0_b_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4629 \$6097 \$7032 \$7106 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4630 \$7107 \$7032 \$6098 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4631 b6_r0_b \$7034 \$7107 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4632 \$6097 \$7033 b6_r0_b vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P
+ AD=0.2562P PS=2.06U PD=2.06U
M$4633 \$7267
+ b7_not|b7_q0_not|b7_q1_not|b7_q2_not|b7_q3_not|b7_q4_not|b7_q5_not|b7_q6_not|b7_q7_not
+ \$6957 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4634 \$7264 a0|b0_p0|b1_p0|b2_p0|b3_p0|b4_p0|b5_p0|b6_p0|b7_p0 \$7267 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4635 \$6959 b1_q3|b7|b7_q0|b7_q1|b7_q2|b7_q4|b7_q5|b7_q6|b7_q7 \$7264 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4636 \$7265 b1_q3|b7|b7_q0|b7_q1|b7_q2|b7_q4|b7_q5|b7_q6|b7_q7 \$6957 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4637 \$6958 a0|b0_p0|b1_p0|b2_p0|b3_p0|b4_p0|b5_p0|b6_p0|b7_p0 \$7265 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4638 \$6959
+ b7_not|b7_q0_not|b7_q1_not|b7_q2_not|b7_q3_not|b7_q4_not|b7_q5_not|b7_q6_not|b7_q7_not
+ \$6958 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4639 \$6211 \$7040 \$7267 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4640 \$7109 \$7041 \$6211 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4641 \$6958 \$7039 \$7109 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4642 \$7110 \$7039 \$7267 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4643 \$6427 \$7041 \$7110 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4644 \$6958 \$7040 \$6427 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4645 \$6960 \$7040 \$6105 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4646 \$7111 \$7041 \$6960 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4647 \$6104 \$7039 \$7111 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4648 \$7112 \$7039 \$6105 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4649 \$6961 \$7041 \$7112 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4650 \$6104 \$7040 \$6961 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P
+ PS=2.06U PD=2.06U
M$4651 p0_not
+ a0_not|b0_p0_not|b1_p0_not|b2_p0_not|b3_p0_not|b5_p0_not|b6_p0_not|b7_p0_not
+ b0_c0_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$4652 p0_not
+ b0_not|b0_q0_not|b0_q1_not|b0_q3_not|b0_q4_not|b0_q5_not|b0_q6_not|b0_q7_not|b1_q2_not
+ b0_c0_not vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U
+ PD=2.06U
M$4653 \$7737 a0|b0_p0|b1_p0|b2_p0|b3_p0|b4_p0|b5_p0|b6_p0|b7_p0 p0_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4654 b0_c0 b0|b0_q0|b0_q1|b0_q2|b0_q3|b0_q4|b0_q5|b0_q6|b0_q7 \$7737 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4655 \$7739 b0|b0_q0|b0_q1|b0_q2|b0_q3|b0_q4|b0_q5|b0_q6|b0_q7 b0_c0_not vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4656 p0 a0|b0_p0|b1_p0|b2_p0|b3_p0|b4_p0|b5_p0|b6_p0|b7_p0 \$7739 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4657 b0_c0
+ b0_not|b0_q0_not|b0_q1_not|b0_q3_not|b0_q4_not|b0_q5_not|b0_q6_not|b0_q7_not|b1_q2_not
+ p0 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4658 b0_c0
+ a0_not|b0_p0_not|b1_p0_not|b2_p0_not|b3_p0_not|b5_p0_not|b6_p0_not|b7_p0_not
+ p0 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4659 \$7254
+ b5_not|b5_q0_not|b5_q1_not|b5_q2_not|b5_q3_not|b5_q4_not|b5_q5_not|b5_q6_not|b5_q7_not
+ \$6948 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4660 \$7251 a0|b0_p0|b1_p0|b2_p0|b3_p0|b4_p0|b5_p0|b6_p0|b7_p0 \$7254 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4661 \$6950 b5|b5_q0|b5_q1|b5_q2|b5_q3|b5_q4|b5_q5|b5_q6|b5_q7 \$7251 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4662 \$7252 b5|b5_q0|b5_q1|b5_q2|b5_q3|b5_q4|b5_q5|b5_q6|b5_q7 \$6948 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4663 \$6949 a0|b0_p0|b1_p0|b2_p0|b3_p0|b4_p0|b5_p0|b6_p0|b7_p0 \$7252 vss
+ nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
M$4664 \$6950
+ b5_not|b5_q0_not|b5_q1_not|b5_q2_not|b5_q3_not|b5_q4_not|b5_q5_not|b5_q6_not|b5_q7_not
+ \$6949 vss nfet_03v3 L=0.28U W=0.42U AS=0.2562P AD=0.2562P PS=2.06U PD=2.06U
.ENDS 8b_mult
