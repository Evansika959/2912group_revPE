VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fa8b_rev
  CLASS BLOCK ;
  FOREIGN fa8b_rev ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.665 BY 212.100 ;
  PIN c_8_not
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 104.010 24.915 108.095 25.250 ;
    END
  END c_8_not
  PIN z
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 100.280 27.290 111.325 27.590 ;
    END
  END z
  PIN z_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT 102.630 26.755 108.680 27.025 ;
    END
  END z_not
  PIN c0
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 161.170 184.800 164.390 185.100 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 30.005 181.695 50.350 181.990 ;
    END
  END c0
  PIN c0_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 158.225 184.055 165.950 184.355 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 29.825 180.830 50.935 181.125 ;
    END
  END c0_not
  PIN s0
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 152.405 180.965 162.485 181.300 ;
    END
  END s0
  PIN s0_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 159.755 183.040 162.485 183.315 ;
    END
  END s0_not
  PIN s1
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 152.205 161.240 162.285 161.575 ;
    END
  END s1
  PIN s1_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 159.555 163.315 162.285 163.590 ;
    END
  END s1_not
  PIN s2
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 152.360 141.595 162.440 141.930 ;
    END
  END s2
  PIN s2_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 159.710 143.670 162.440 143.945 ;
    END
  END s2_not
  PIN s3
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 152.360 121.800 162.440 122.135 ;
    END
  END s3
  PIN s3_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 159.710 123.875 162.440 124.150 ;
    END
  END s3_not
  PIN s4
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 152.280 102.045 162.360 102.380 ;
    END
  END s4
  PIN s4_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 159.630 104.120 162.360 104.395 ;
    END
  END s4_not
  PIN s5
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 152.385 82.330 162.465 82.665 ;
    END
  END s5
  PIN s5_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 159.735 84.405 162.465 84.680 ;
    END
  END s5_not
  PIN s6
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 152.385 62.360 162.465 62.695 ;
    END
  END s6
  PIN s6_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 159.735 64.435 162.465 64.710 ;
    END
  END s6_not
  PIN s7
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 152.385 42.695 162.465 43.030 ;
    END
  END s7
  PIN s7_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 159.735 44.770 162.465 45.045 ;
    END
  END s7_not
  PIN VDD
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 25.150 190.475 105.170 191.390 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 25.035 170.700 105.185 171.615 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 25.070 151.075 105.170 151.990 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 25.045 131.270 105.185 132.185 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 24.985 111.465 105.195 112.380 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 25.030 91.800 105.145 92.715 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 25.070 71.830 105.170 72.745 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 25.015 52.165 105.200 53.080 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 25.000 34.230 105.215 35.475 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 105.495 34.230 170.195 35.475 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 105.480 52.165 170.210 53.080 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 105.450 71.830 170.265 72.745 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 105.425 91.800 170.225 92.715 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 105.475 111.465 170.180 112.380 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 105.465 131.270 170.240 132.185 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 105.450 151.075 170.265 151.990 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 105.465 170.700 170.230 171.615 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 105.450 190.475 170.345 191.390 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 25.025 175.390 95.930 176.305 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 25.060 155.675 95.905 156.590 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 25.045 136.050 95.945 136.965 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 26.610 115.835 26.620 115.845 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 24.995 96.470 95.860 97.385 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 25.015 76.750 95.835 77.665 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 25.050 56.810 96.010 57.725 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 24.965 37.140 95.970 38.040 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 25.000 19.160 95.920 20.405 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 96.210 175.390 170.220 176.305 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 96.185 155.675 170.255 156.590 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 96.225 136.050 170.240 136.965 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 96.155 116.245 170.175 117.160 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 96.140 96.470 170.190 97.385 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 96.115 76.750 170.210 77.665 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 96.290 56.810 170.245 57.725 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 96.250 37.140 170.145 38.040 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 96.200 19.160 170.180 20.405 ;
    END
  END VSS
  PIN c_8
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal3 ;
        RECT 118.430 18.370 119.455 18.720 ;
    END
  END c_8
  PIN a0_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 32.960 184.850 35.420 185.155 ;
    END
  END a0_f
  PIN a0_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 32.920 184.115 35.425 184.410 ;
    END
  END a0_not_f
  PIN a0_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 146.970 189.670 162.705 190.080 ;
    END
  END a0_b
  PIN a0_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 147.565 188.890 162.695 189.345 ;
    END
  END a0_not_b
  PIN a7_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 32.830 46.535 35.290 46.840 ;
    END
  END a7_f
  PIN a7_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 32.790 45.800 35.295 46.095 ;
    END
  END a7_not_f
  PIN a7_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 146.950 51.400 162.685 51.810 ;
    END
  END a7_b
  PIN a7_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 147.545 50.620 162.675 51.075 ;
    END
  END a7_not_b
  PIN b0
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 32.925 183.400 35.440 183.695 ;
    END
  END b0
  PIN b0_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 32.960 182.770 35.425 183.065 ;
    END
  END b0_not
  PIN a1
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 32.915 165.160 35.375 165.465 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 146.770 169.945 162.505 170.355 ;
    END
  END a1
  PIN a1_not
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 32.875 164.425 35.380 164.720 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 147.365 169.165 162.495 169.620 ;
    END
  END a1_not
  PIN b1
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 32.880 163.710 35.395 164.005 ;
    END
  END b1
  PIN b1_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 32.915 163.080 35.380 163.375 ;
    END
  END b1_not
  PIN a2
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 33.105 145.450 35.565 145.755 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 146.925 150.300 162.660 150.710 ;
    END
  END a2
  PIN a2_not
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 33.065 144.715 35.570 145.010 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 147.520 149.520 162.650 149.975 ;
    END
  END a2_not
  PIN b2
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 33.070 144.000 35.585 144.295 ;
    END
  END b2
  PIN b2_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 33.105 143.370 35.570 143.665 ;
    END
  END b2_not
  PIN a3
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 32.910 125.610 35.370 125.915 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 146.925 130.505 162.660 130.915 ;
    END
  END a3
  PIN a3_not
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 32.870 124.875 35.375 125.170 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 147.520 129.725 162.650 130.180 ;
    END
  END a3_not
  PIN b3
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 32.875 124.160 35.390 124.455 ;
    END
  END b3
  PIN b3_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 32.910 123.530 35.375 123.825 ;
    END
  END b3_not
  PIN a4
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 32.780 105.900 35.240 106.205 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 146.845 110.750 162.580 111.160 ;
    END
  END a4
  PIN a4_not
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 32.740 105.165 35.245 105.460 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 147.440 109.970 162.570 110.425 ;
    END
  END a4_not
  PIN b4
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 32.745 104.450 35.260 104.745 ;
    END
  END b4
  PIN b4_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 32.780 103.820 35.245 104.115 ;
    END
  END b4_not
  PIN a5
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 32.910 86.140 35.370 86.445 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 146.950 91.035 162.685 91.445 ;
    END
  END a5
  PIN a5_not
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 32.870 85.405 35.375 85.700 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 147.545 90.255 162.675 90.710 ;
    END
  END a5_not
  PIN b5
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 32.875 84.690 35.390 84.985 ;
    END
  END b5
  PIN b5_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 32.910 84.060 35.375 84.355 ;
    END
  END b5_not
  PIN a6
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 32.860 66.330 35.320 66.635 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 146.950 71.065 162.685 71.475 ;
    END
  END a6
  PIN a6_not
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 32.820 65.595 35.325 65.890 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 147.545 70.285 162.675 70.740 ;
    END
  END a6_not
  PIN b6
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 32.825 64.880 35.340 65.175 ;
    END
  END b6
  PIN b6_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 32.860 64.250 35.325 64.545 ;
    END
  END b6_not
  PIN b7
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 32.795 45.085 35.310 45.380 ;
    END
  END b7
  PIN b7_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 32.830 44.455 35.295 44.750 ;
    END
  END b7_not
  OBS
      LAYER Nwell ;
        RECT 33.240 19.365 162.485 191.395 ;
      LAYER Metal1 ;
        RECT 33.670 185.400 165.930 191.395 ;
        RECT 33.670 184.655 160.870 185.400 ;
        RECT 164.690 184.655 165.930 185.400 ;
        RECT 33.670 183.755 157.925 184.655 ;
        RECT 33.670 183.615 165.930 183.755 ;
        RECT 33.670 182.740 159.455 183.615 ;
        RECT 162.785 182.740 165.930 183.615 ;
        RECT 33.670 181.600 165.930 182.740 ;
        RECT 33.670 180.665 152.105 181.600 ;
        RECT 162.785 180.665 165.930 181.600 ;
        RECT 33.670 163.890 165.930 180.665 ;
        RECT 33.670 163.015 159.255 163.890 ;
        RECT 162.585 163.015 165.930 163.890 ;
        RECT 33.670 161.875 165.930 163.015 ;
        RECT 33.670 160.940 151.905 161.875 ;
        RECT 162.585 160.940 165.930 161.875 ;
        RECT 33.670 144.245 165.930 160.940 ;
        RECT 33.670 143.370 159.410 144.245 ;
        RECT 162.740 143.370 165.930 144.245 ;
        RECT 33.670 142.230 165.930 143.370 ;
        RECT 33.670 141.295 152.060 142.230 ;
        RECT 162.740 141.295 165.930 142.230 ;
        RECT 33.670 124.450 165.930 141.295 ;
        RECT 33.670 123.575 159.410 124.450 ;
        RECT 162.740 123.575 165.930 124.450 ;
        RECT 33.670 122.435 165.930 123.575 ;
        RECT 33.670 121.500 152.060 122.435 ;
        RECT 162.740 121.500 165.930 122.435 ;
        RECT 33.670 104.695 165.930 121.500 ;
        RECT 33.670 103.820 159.330 104.695 ;
        RECT 162.660 103.820 165.930 104.695 ;
        RECT 33.670 102.680 165.930 103.820 ;
        RECT 33.670 101.745 151.980 102.680 ;
        RECT 162.660 101.745 165.930 102.680 ;
        RECT 33.670 84.980 165.930 101.745 ;
        RECT 33.670 84.105 159.435 84.980 ;
        RECT 162.765 84.105 165.930 84.980 ;
        RECT 33.670 82.965 165.930 84.105 ;
        RECT 33.670 82.030 152.085 82.965 ;
        RECT 162.765 82.030 165.930 82.965 ;
        RECT 33.670 65.010 165.930 82.030 ;
        RECT 33.670 64.135 159.435 65.010 ;
        RECT 162.765 64.135 165.930 65.010 ;
        RECT 33.670 62.995 165.930 64.135 ;
        RECT 33.670 62.060 152.085 62.995 ;
        RECT 162.765 62.060 165.930 62.995 ;
        RECT 33.670 45.345 165.930 62.060 ;
        RECT 33.670 44.470 159.435 45.345 ;
        RECT 162.765 44.470 165.930 45.345 ;
        RECT 33.670 43.330 165.930 44.470 ;
        RECT 33.670 42.395 152.085 43.330 ;
        RECT 162.765 42.395 165.930 43.330 ;
        RECT 33.670 27.890 165.930 42.395 ;
        RECT 33.670 26.990 99.980 27.890 ;
        RECT 111.625 26.990 165.930 27.890 ;
        RECT 33.670 26.455 102.330 26.990 ;
        RECT 108.980 26.455 165.930 26.990 ;
        RECT 33.670 25.550 165.930 26.455 ;
        RECT 33.670 24.615 103.710 25.550 ;
        RECT 108.395 24.615 165.930 25.550 ;
        RECT 33.670 19.360 165.930 24.615 ;
      LAYER Metal2 ;
        RECT 29.910 18.290 165.840 191.395 ;
      LAYER Metal3 ;
        RECT 24.980 189.370 146.670 190.175 ;
        RECT 163.005 189.370 166.555 190.175 ;
        RECT 24.980 188.590 147.265 189.370 ;
        RECT 162.995 188.590 166.555 189.370 ;
        RECT 24.980 185.455 166.555 188.590 ;
        RECT 24.980 184.710 32.660 185.455 ;
        RECT 35.720 184.710 166.555 185.455 ;
        RECT 24.980 183.815 32.620 184.710 ;
        RECT 35.725 183.995 166.555 184.710 ;
        RECT 24.980 183.100 32.625 183.815 ;
        RECT 35.740 183.100 166.555 183.995 ;
        RECT 24.980 182.470 32.660 183.100 ;
        RECT 35.725 182.470 166.555 183.100 ;
        RECT 24.980 182.290 166.555 182.470 ;
        RECT 24.980 181.425 29.705 182.290 ;
        RECT 50.650 181.425 166.555 182.290 ;
        RECT 24.980 180.530 29.525 181.425 ;
        RECT 51.235 180.530 166.555 181.425 ;
        RECT 24.980 176.605 166.555 180.530 ;
        RECT 24.980 171.915 166.555 175.090 ;
        RECT 24.980 169.645 146.470 170.400 ;
        RECT 162.805 169.645 166.555 170.400 ;
        RECT 24.980 168.865 147.065 169.645 ;
        RECT 162.795 168.865 166.555 169.645 ;
        RECT 24.980 165.765 166.555 168.865 ;
        RECT 24.980 165.020 32.615 165.765 ;
        RECT 35.675 165.020 166.555 165.765 ;
        RECT 24.980 164.125 32.575 165.020 ;
        RECT 35.680 164.305 166.555 165.020 ;
        RECT 24.980 163.410 32.580 164.125 ;
        RECT 35.695 163.410 166.555 164.305 ;
        RECT 24.980 162.780 32.615 163.410 ;
        RECT 35.680 162.780 166.555 163.410 ;
        RECT 24.980 156.890 166.555 162.780 ;
        RECT 24.980 152.290 166.555 155.375 ;
        RECT 24.980 150.000 146.625 150.775 ;
        RECT 162.960 150.000 166.555 150.775 ;
        RECT 24.980 149.220 147.220 150.000 ;
        RECT 162.950 149.220 166.555 150.000 ;
        RECT 24.980 146.055 166.555 149.220 ;
        RECT 24.980 145.310 32.805 146.055 ;
        RECT 35.865 145.310 166.555 146.055 ;
        RECT 24.980 144.415 32.765 145.310 ;
        RECT 35.870 144.595 166.555 145.310 ;
        RECT 24.980 143.700 32.770 144.415 ;
        RECT 35.885 143.700 166.555 144.595 ;
        RECT 24.980 143.070 32.805 143.700 ;
        RECT 35.870 143.070 166.555 143.700 ;
        RECT 24.980 137.265 166.555 143.070 ;
        RECT 24.980 132.485 166.555 135.750 ;
        RECT 24.980 130.205 146.625 130.970 ;
        RECT 162.960 130.205 166.555 130.970 ;
        RECT 24.980 129.425 147.220 130.205 ;
        RECT 162.950 129.425 166.555 130.205 ;
        RECT 24.980 126.215 166.555 129.425 ;
        RECT 24.980 125.470 32.610 126.215 ;
        RECT 35.670 125.470 166.555 126.215 ;
        RECT 24.980 124.575 32.570 125.470 ;
        RECT 35.675 124.755 166.555 125.470 ;
        RECT 24.980 123.860 32.575 124.575 ;
        RECT 35.690 123.860 166.555 124.755 ;
        RECT 24.980 123.230 32.610 123.860 ;
        RECT 35.675 123.230 166.555 123.860 ;
        RECT 24.980 117.460 166.555 123.230 ;
        RECT 24.980 116.145 95.855 117.460 ;
        RECT 24.980 115.535 26.310 116.145 ;
        RECT 26.920 115.945 95.855 116.145 ;
        RECT 26.920 115.535 166.555 115.945 ;
        RECT 24.980 112.680 166.555 115.535 ;
        RECT 24.980 110.450 146.545 111.165 ;
        RECT 162.880 110.450 166.555 111.165 ;
        RECT 24.980 109.670 147.140 110.450 ;
        RECT 162.870 109.670 166.555 110.450 ;
        RECT 24.980 106.505 166.555 109.670 ;
        RECT 24.980 105.760 32.480 106.505 ;
        RECT 35.540 105.760 166.555 106.505 ;
        RECT 24.980 104.865 32.440 105.760 ;
        RECT 35.545 105.045 166.555 105.760 ;
        RECT 24.980 104.150 32.445 104.865 ;
        RECT 35.560 104.150 166.555 105.045 ;
        RECT 24.980 103.520 32.480 104.150 ;
        RECT 35.545 103.520 166.555 104.150 ;
        RECT 24.980 97.685 166.555 103.520 ;
        RECT 24.980 93.015 166.555 96.170 ;
        RECT 24.980 90.735 146.650 91.500 ;
        RECT 162.985 90.735 166.555 91.500 ;
        RECT 24.980 89.955 147.245 90.735 ;
        RECT 162.975 89.955 166.555 90.735 ;
        RECT 24.980 86.745 166.555 89.955 ;
        RECT 24.980 86.000 32.610 86.745 ;
        RECT 35.670 86.000 166.555 86.745 ;
        RECT 24.980 85.105 32.570 86.000 ;
        RECT 35.675 85.285 166.555 86.000 ;
        RECT 24.980 84.390 32.575 85.105 ;
        RECT 35.690 84.390 166.555 85.285 ;
        RECT 24.980 83.760 32.610 84.390 ;
        RECT 35.675 83.760 166.555 84.390 ;
        RECT 24.980 77.965 166.555 83.760 ;
        RECT 24.980 73.045 166.555 76.450 ;
        RECT 24.980 70.765 146.650 71.530 ;
        RECT 162.985 70.765 166.555 71.530 ;
        RECT 24.980 69.985 147.245 70.765 ;
        RECT 162.975 69.985 166.555 70.765 ;
        RECT 24.980 66.935 166.555 69.985 ;
        RECT 24.980 66.190 32.560 66.935 ;
        RECT 35.620 66.190 166.555 66.935 ;
        RECT 24.980 65.295 32.520 66.190 ;
        RECT 35.625 65.475 166.555 66.190 ;
        RECT 24.980 64.580 32.525 65.295 ;
        RECT 35.640 64.580 166.555 65.475 ;
        RECT 24.980 63.950 32.560 64.580 ;
        RECT 35.625 63.950 166.555 64.580 ;
        RECT 24.980 58.025 166.555 63.950 ;
        RECT 24.980 53.380 166.555 56.510 ;
        RECT 24.980 51.100 146.650 51.865 ;
        RECT 162.985 51.100 166.555 51.865 ;
        RECT 24.980 50.320 147.245 51.100 ;
        RECT 162.975 50.320 166.555 51.100 ;
        RECT 24.980 47.140 166.555 50.320 ;
        RECT 24.980 46.395 32.530 47.140 ;
        RECT 35.590 46.395 166.555 47.140 ;
        RECT 24.980 45.500 32.490 46.395 ;
        RECT 35.595 45.680 166.555 46.395 ;
        RECT 24.980 44.785 32.495 45.500 ;
        RECT 35.610 44.785 166.555 45.680 ;
        RECT 24.980 44.155 32.530 44.785 ;
        RECT 35.595 44.155 166.555 44.785 ;
        RECT 24.980 38.340 166.555 44.155 ;
        RECT 24.980 35.775 166.555 36.840 ;
        RECT 24.980 20.705 166.555 33.930 ;
        RECT 24.980 18.370 118.130 18.860 ;
        RECT 119.755 18.370 166.555 18.860 ;
  END
END fa8b_rev
END LIBRARY

