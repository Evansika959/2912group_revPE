`default_nettype none

module fa16_rev_wrapped (
    `ifdef USE_POWER_PINS
    inout wire vdd,
    inout wire vss,
    `endif

    // Input ports
    inout  wire [15:0] a,
    inout  wire [15:0] a_not,
    inout  wire [15:0] b,
    inout  wire [15:0] b_not,
    inout  wire        c0_f,
    inout  wire        c0_f_not,
    inout  wire        c15,
    inout  wire        c15_not,

    // Output ports
    inout wire [15:0] s,
    inout wire [15:0] s_not,
    inout wire [15:0] a_b,
    inout wire [15:0] a_not_b,
    inout wire        z,
    inout wire        z_not,
    inout wire        c0_b,
    inout wire        c0_not_b,
);

    // Power handling
    `ifndef USE_POWER_PINS
    wire vdd = 1'b1;
    wire vss = 1'b0;
    `endif

    // Unused macro pins preserved to track full LEF interface
    wire unused_z;
    wire unused_z_not;
    wire unused_c0_b;
    wire unused_c0_not_b;

    (* keep *)
    fa16b_rev u_fa16b_rev (
        .z           (unused_z),
        .z_not       (unused_z_not),
        .c0_b        (unused_c0_b),
        .c0_not_b    (unused_c0_not_b),
        .c15_not     (c15_not),
        .c15         (c15),
        .s5_not      (s_not[5]),
        .s5          (s[5]),
        .s0_not      (s_not[0]),
        .s0          (s[0]),
        .s6_not      (s_not[6]),
        .s6          (s[6]),
        .s1_not      (s_not[1]),
        .s1          (s[1]),
        .s7_not      (s_not[7]),
        .s7          (s[7]),
        .s2_not      (s_not[2]),
        .s2          (s[2]),
        .s8_not      (s_not[8]),
        .s8          (s[8]),
        .s3_not      (s_not[3]),
        .s3          (s[3]),
        .s9_not      (s_not[9]),
        .s9          (s[9]),
        .s4_not      (s_not[4]),
        .s4          (s[4]),
        .s10_not     (s_not[10]),
        .s10         (s[10]),
        .s11_not     (s_not[11]),
        .s11         (s[11]),
        .s12_not     (s_not[12]),
        .s12         (s[12]),
        .s13_not     (s_not[13]),
        .s13         (s[13]),
        .s14_not     (s_not[14]),
        .s14         (s[14]),
        .s15_not     (s_not[15]),
        .s15         (s[15]),
        .c0_f        (c0_f),
        .c0_f_not    (c0_f_not),
        .vss         (vss),
        .vdd         (vdd),
        .a0_f        (a[0]),
        .a0_not_f    (a_not[0]),
        .b0          (b[0]),
        .b0_not      (b_not[0]),
        .a1_f        (a[1]),
        .a1_not_f    (a_not[1]),
        .b1          (b[1]),
        .b1_not      (b_not[1]),
        .a2_f        (a[2]),
        .a2_not_f    (a_not[2]),
        .b2          (b[2]),
        .b2_not      (b_not[2]),
        .a3_f        (a[3]),
        .a3_not_f    (a_not[3]),
        .b3          (b[3]),
        .b3_not      (b_not[3]),
        .a4_f        (a[4]),
        .a4_not_f    (a_not[4]),
        .b4          (b[4]),
        .b4_not      (b_not[4]),
        .a5_f        (a[5]),
        .a5_not_f    (a_not[5]),
        .b5          (b[5]),
        .b5_not      (b_not[5]),
        .a6_f        (a[6]),
        .a6_not_f    (a_not[6]),
        .b6          (b[6]),
        .b6_not      (b_not[6]),
        .a7_f        (a[7]),
        .a7_not_f    (a_not[7]),
        .b7          (b[7]),
        .b7_not      (b_not[7]),
        .a8_f        (a[8]),
        .a8_not_f    (a_not[8]),
        .b8          (b[8]),
        .b8_not      (b_not[8]),
        .a9_f        (a[9]),
        .a9_not_f    (a_not[9]),
        .b9          (b[9]),
        .b9_not      (b_not[9]),
        .a10_f       (a[10]),
        .a10_not_f   (a_not[10]),
        .b10         (b[10]),
        .b10_not     (b_not[10]),
        .a11_f       (a[11]),
        .a11_not_f   (a_not[11]),
        .b11         (b[11]),
        .b11_not     (b_not[11]),
        .a12_f       (a[12]),
        .a12_not_f   (a_not[12]),
        .b12         (b[12]),
        .b12_not     (b_not[12]),
        .a13_f       (a[13]),
        .a13_not_f   (a_not[13]),
        .b13         (b[13]),
        .b13_not     (b_not[13]),
        .a14_f       (a[14]),
        .a14_not_f   (a_not[14]),
        .b14         (b[14]),
        .b14_not     (b_not[14]),
        .a15_f       (a[15]),
        .a15_not_f   (a_not[15]),
        .b15         (b[15]),
        .b15_not     (b_not[15]),
        .a0_b        (a_b[0]),
        .a0_not_b    (a_not_b[0]),
        .a1_b        (a_b[1]),
        .a1_not_b    (a_not_b[1]),
        .a2_b        (a_b[2]),
        .a2_not_b    (a_not_b[2]),
        .a3_b        (a_b[3]),
        .a3_not_b    (a_not_b[3]),
        .a4_b        (a_b[4]),
        .a4_not_b    (a_not_b[4]),
        .a5_b        (a_b[5]),
        .a5_not_b    (a_not_b[5]),
        .a6_b        (a_b[6]),
        .a6_not_b    (a_not_b[6]),
        .a7_b        (a_b[7]),
        .a7_not_b    (a_not_b[7]),
        .a8_b        (a_b[8]),
        .a8_not_b    (a_not_b[8]),
        .a9_b        (a_b[9]),
        .a9_not_b    (a_not_b[9]),
        .a10_b       (a_b[10]),
        .a10_not_b   (a_not_b[10]),
        .a11_b       (a_b[11]),
        .a11_not_b   (a_not_b[11]),
        .a12_b       (a_b[12]),
        .a12_not_b   (a_not_b[12]),
        .a13_b       (a_b[13]),
        .a13_not_b   (a_not_b[13]),
        .a14_b       (a_b[14]),
        .a14_not_b   (a_not_b[14]),
        .a15_b       (a_b[15]),
        .a15_not_b   (a_not_b[15])
    );

endmodule