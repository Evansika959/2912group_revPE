* NGSPICE file created from 16b_FA.ext - technology: gf180mcuD

.subckt pfet$1 a_28_144# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_144# a_n92_0# w_n180_n88# pfet_03v3 ad=0.273p pd=2.14u as=0.273p ps=2.14u w=0.42u l=0.28u
.ends

.subckt nfet$1$1 a_n84_0# a_94_0# a_30_144# VSUBS
X0 a_94_0# a_30_144# a_n84_0# VSUBS nfet_03v3 ad=0.2562p pd=2.06u as=0.2562p ps=2.06u w=0.42u l=0.28u
.ends

.subckt MAJ w_26_1560# a_551_708# a_7235_2410# a_4594_2030# a_3643_708# a_11429_1029#
+ a_639_1698# a_2043_2038# a_644_83# m1_7413_2589# a_5135_2038# a_1502_2030# pfet$1_7/VSUBS
+ a_749_2028#
Xpfet$1_6 a_7235_2410# w_26_1560# a_644_83# a_11429_1029# pfet$1
Xnfet$1$1_1 m1_10043_1029# a_639_1698# a_749_2028# pfet$1_7/VSUBS nfet$1$1
Xpfet$1_7 a_7235_2410# w_26_1560# m1_7413_2589# a_639_1698# pfet$1
Xnfet$1$1_2 a_644_83# a_11429_1029# a_2043_2038# pfet$1_7/VSUBS nfet$1$1
Xnfet$1$1_3 m1_8218_1029# m1_7413_2589# a_7235_2410# pfet$1_7/VSUBS nfet$1$1
Xnfet$1$1_4 a_11429_1029# m1_10043_1029# a_7235_2410# pfet$1_7/VSUBS nfet$1$1
Xnfet$1$1_5 a_644_83# m1_8218_1029# a_749_2028# pfet$1_7/VSUBS nfet$1$1
Xnfet$1$1_6 a_644_83# a_11429_1029# a_5135_2038# pfet$1_7/VSUBS nfet$1$1
Xnfet$1$1_7 m1_7413_2589# a_639_1698# a_2043_2038# pfet$1_7/VSUBS nfet$1$1
Xpfet$1_0 a_749_2028# w_26_1560# m1_7413_2589# a_639_1698# pfet$1
Xpfet$1_1 a_2043_2038# w_26_1560# m1_8223_2129# m1_7413_2589# pfet$1
Xpfet$1_3 a_5135_2038# w_26_1560# m1_10121_2129# a_639_1698# pfet$1
Xpfet$1_2 a_5135_2038# w_26_1560# a_644_83# m1_8223_2129# pfet$1
Xpfet$1_4 a_2043_2038# w_26_1560# a_11429_1029# m1_10121_2129# pfet$1
Xpfet$1_5 a_749_2028# w_26_1560# a_644_83# a_11429_1029# pfet$1
Xnfet$1$1_0 m1_7413_2589# a_639_1698# a_5135_2038# pfet$1_7/VSUBS nfet$1$1
X0 a_2043_2038# a_644_83# a_1502_2030# pfet$1_7/VSUBS nfet_03v3 ad=0.64155p pd=3.67u as=0.64837p ps=3.68u w=1.365u l=0.55u
X1 a_3643_708# a_639_1698# a_5135_2038# pfet$1_7/VSUBS nfet_03v3 ad=0.6925p pd=3.77u as=0.67172p ps=3.74u w=1.385u l=0.55u
X2 a_4594_2030# a_644_83# a_7235_2410# w_26_1560# pfet_03v3 ad=0.60515p pd=3.45u as=0.6669p ps=3.55u w=1.235u l=0.5u
X3 a_7235_2410# a_644_83# a_3643_708# pfet$1_7/VSUBS nfet_03v3 ad=0.6576p pd=3.7u as=0.63705p ps=3.67u w=1.37u l=0.55u
X4 a_749_2028# a_644_83# a_551_708# pfet$1_7/VSUBS nfet_03v3 ad=0.6576p pd=3.7u as=0.63705p ps=3.67u w=1.37u l=0.55u
X5 a_5135_2038# a_639_1698# a_4594_2030# w_26_1560# pfet_03v3 ad=0.60515p pd=3.45u as=0.64837p ps=3.52u w=1.235u l=0.5u
X6 a_5135_2038# a_644_83# a_4594_2030# pfet$1_7/VSUBS nfet_03v3 ad=0.64155p pd=3.67u as=0.64837p ps=3.68u w=1.365u l=0.55u
X7 a_1502_2030# a_639_1698# a_749_2028# pfet$1_7/VSUBS nfet_03v3 ad=0.65797p pd=3.76u as=0.74287p ps=3.88u w=1.415u l=0.55u
X8 a_551_708# a_639_1698# a_2043_2038# pfet$1_7/VSUBS nfet_03v3 ad=0.6925p pd=3.77u as=0.67172p ps=3.74u w=1.385u l=0.55u
X9 a_1502_2030# a_644_83# a_749_2028# w_26_1560# pfet_03v3 ad=0.60515p pd=3.45u as=0.6669p ps=3.55u w=1.235u l=0.5u
X10 a_551_708# a_644_83# a_2043_2038# w_26_1560# pfet_03v3 ad=0.70395p pd=3.61u as=0.6422p ps=3.51u w=1.235u l=0.5u
X11 a_749_2028# a_639_1698# a_551_708# w_26_1560# pfet_03v3 ad=0.6669p pd=3.55u as=0.60515p ps=3.45u w=1.235u l=0.5u
X12 a_2043_2038# a_639_1698# a_1502_2030# w_26_1560# pfet_03v3 ad=0.60515p pd=3.45u as=0.64837p ps=3.52u w=1.235u l=0.5u
X13 a_7235_2410# a_639_1698# a_3643_708# w_26_1560# pfet_03v3 ad=0.6669p pd=3.55u as=0.60515p ps=3.45u w=1.235u l=0.5u
X14 a_4594_2030# a_639_1698# a_7235_2410# pfet$1_7/VSUBS nfet_03v3 ad=0.65797p pd=3.76u as=0.74287p ps=3.88u w=1.415u l=0.55u
X15 a_3643_708# a_644_83# a_5135_2038# w_26_1560# pfet_03v3 ad=0.70395p pd=3.61u as=0.6422p ps=3.51u w=1.235u l=0.5u
.ends

.subckt pfet a_28_144# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_144# a_n92_0# w_n180_n88# pfet_03v3 ad=0.273p pd=2.14u as=0.273p ps=2.14u w=0.42u l=0.28u
.ends

.subckt nfet$1 a_n84_0# a_94_0# a_30_144# VSUBS
X0 a_94_0# a_30_144# a_n84_0# VSUBS nfet_03v3 ad=0.2562p pd=2.06u as=0.2562p ps=2.06u w=0.42u l=0.28u
.ends

.subckt UMA a_319_1607# a_4705_1617# a_209_1277# a_3411_1607# a_n806_2017# a_n690_608#
+ pfet_7/VSUBS a_121_287# m1_n6688_1443# a_1613_1617# a_3213_287# w_n5735_1139# a_4164_1609#
+ a_n912_608#
Xpfet_0 a_4164_1609# w_n5735_1139# a_209_1277# m1_n6688_1443# pfet
Xpfet_1 a_3213_287# w_n5735_1139# m1_n4118_1708# a_209_1277# pfet
Xpfet_2 a_121_287# w_n5735_1139# a_n690_608# m1_n4118_1708# pfet
Xpfet_4 a_3213_287# w_n5735_1139# a_n912_608# m1_n2220_1708# pfet
Xpfet_3 a_121_287# w_n5735_1139# m1_n2220_1708# m1_n6688_1443# pfet
Xpfet_5 a_4164_1609# w_n5735_1139# a_n690_608# a_n912_608# pfet
Xpfet_6 a_n806_2017# w_n5735_1139# a_n690_608# a_n912_608# pfet
Xpfet_7 a_n806_2017# w_n5735_1139# a_209_1277# m1_n6688_1443# pfet
Xnfet$1_0 a_209_1277# m1_n6688_1443# a_121_287# pfet_7/VSUBS nfet$1
Xnfet$1_1 m1_n2298_608# m1_n6688_1443# a_4164_1609# pfet_7/VSUBS nfet$1
Xnfet$1_2 a_n690_608# a_n912_608# a_3213_287# pfet_7/VSUBS nfet$1
Xnfet$1_3 m1_n4123_608# a_209_1277# a_n806_2017# pfet_7/VSUBS nfet$1
Xnfet$1_4 a_n912_608# m1_n2298_608# a_n806_2017# pfet_7/VSUBS nfet$1
Xnfet$1_5 a_n690_608# m1_n4123_608# a_4164_1609# pfet_7/VSUBS nfet$1
Xnfet$1_6 a_n690_608# a_n912_608# a_121_287# pfet_7/VSUBS nfet$1
Xnfet$1_7 a_209_1277# m1_n6688_1443# a_3213_287# pfet_7/VSUBS nfet$1
X0 a_n806_2017# a_n912_608# a_319_1607# w_n5735_1139# pfet_03v3 ad=0.60515p pd=3.45u as=0.6669p ps=3.55u w=1.235u l=0.5u
X1 a_121_287# a_n912_608# a_1613_1617# w_n5735_1139# pfet_03v3 ad=0.70395p pd=3.61u as=0.6422p ps=3.51u w=1.235u l=0.5u
X2 a_n806_2017# a_209_1277# a_319_1607# pfet_7/VSUBS nfet_03v3 ad=0.65797p pd=3.76u as=0.74287p ps=3.88u w=1.415u l=0.55u
X3 a_319_1607# a_209_1277# a_121_287# w_n5735_1139# pfet_03v3 ad=0.6669p pd=3.55u as=0.60515p ps=3.45u w=1.235u l=0.5u
X4 a_319_1607# a_n912_608# a_121_287# pfet_7/VSUBS nfet_03v3 ad=0.6576p pd=3.7u as=0.63705p ps=3.67u w=1.37u l=0.55u
X5 a_1613_1617# a_209_1277# a_n806_2017# w_n5735_1139# pfet_03v3 ad=0.60515p pd=3.45u as=0.64837p ps=3.52u w=1.235u l=0.5u
X6 a_3411_1607# a_1613_1617# a_3213_287# w_n5735_1139# pfet_03v3 ad=0.6669p pd=3.55u as=0.60515p ps=3.45u w=1.235u l=0.5u
X7 a_4164_1609# a_319_1607# a_3411_1607# w_n5735_1139# pfet_03v3 ad=0.60515p pd=3.45u as=0.6669p ps=3.55u w=1.235u l=0.5u
X8 a_3213_287# a_319_1607# a_4705_1617# w_n5735_1139# pfet_03v3 ad=0.70395p pd=3.61u as=0.6422p ps=3.51u w=1.235u l=0.5u
X9 a_4705_1617# a_1613_1617# a_4164_1609# w_n5735_1139# pfet_03v3 ad=0.60515p pd=3.45u as=0.64837p ps=3.52u w=1.235u l=0.5u
X10 a_121_287# a_209_1277# a_1613_1617# pfet_7/VSUBS nfet_03v3 ad=0.6925p pd=3.77u as=0.67172p ps=3.74u w=1.385u l=0.55u
X11 a_4705_1617# a_319_1607# a_4164_1609# pfet_7/VSUBS nfet_03v3 ad=0.64155p pd=3.67u as=0.64837p ps=3.68u w=1.365u l=0.55u
X12 a_4164_1609# a_1613_1617# a_3411_1607# pfet_7/VSUBS nfet_03v3 ad=0.65797p pd=3.76u as=0.74287p ps=3.88u w=1.415u l=0.55u
X13 a_1613_1617# a_n912_608# a_n806_2017# pfet_7/VSUBS nfet_03v3 ad=0.64155p pd=3.67u as=0.64837p ps=3.68u w=1.365u l=0.55u
X14 a_3213_287# a_1613_1617# a_4705_1617# pfet_7/VSUBS nfet_03v3 ad=0.6925p pd=3.77u as=0.67172p ps=3.74u w=1.385u l=0.55u
X15 a_3411_1607# a_319_1607# a_3213_287# pfet_7/VSUBS nfet_03v3 ad=0.6576p pd=3.7u as=0.63705p ps=3.67u w=1.37u l=0.55u
.ends

.subckt x8b_FA MAJ_7/a_551_708# UMA_7/a_1613_1617# UMA_4/a_4705_1617# MAJ_7/a_1502_2030#
+ MAJ_2/a_1502_2030# UMA_4/a_3411_1607# UMA_0/a_n690_608# MAJ_6/a_644_83# MAJ_2/a_644_83#
+ UMA_0/m1_n6688_1443# UMA_3/a_4705_1617# MAJ_6/a_1502_2030# MAJ_1/a_1502_2030# UMA_0/a_n912_608#
+ MAJ_7/a_3643_708# MAJ_0/m1_7413_2589# UMA_1/a_n912_608# UMA_3/a_3411_1607# MAJ_0/a_639_1698#
+ UMA_2/a_n912_608# MAJ_0/w_26_1560# MAJ_1/a_639_1698# UMA_3/a_n912_608# MAJ_2/a_639_1698#
+ UMA_4/a_n912_608# MAJ_0/a_551_708# MAJ_3/a_639_1698# UMA_5/a_n912_608# UMA_0/a_209_1277#
+ MAJ_7/a_644_83# MAJ_4/a_639_1698# MAJ_7/a_4594_2030# UMA_6/a_n912_608# MAJ_1/w_26_1560#
+ UMA_1/a_209_1277# MAJ_5/a_639_1698# UMA_7/a_4705_1617# UMA_7/a_n912_608# MAJ_3/a_644_83#
+ UMA_2/a_4705_1617# MAJ_6/a_639_1698# UMA_2/a_209_1277# MAJ_5/a_1502_2030# MAJ_1/a_551_708#
+ MAJ_0/a_1502_2030# MAJ_7/a_639_1698# UMA_7/a_319_1607# UMA_3/a_209_1277# UMA_7/a_3411_1607#
+ UMA_4/a_209_1277# MAJ_2/w_26_1560# UMA_2/a_3411_1607# UMA_5/a_209_1277# UMA_6/a_209_1277#
+ MAJ_2/a_551_708# UMA_7/a_209_1277# MAJ_3/w_26_1560# UMA_6/a_4705_1617# UMA_1/a_4705_1617#
+ MAJ_3/a_551_708# MAJ_4/a_1502_2030# MAJ_4/a_644_83# MAJ_4/w_26_1560# MAJ_0/a_11429_1029#
+ UMA_6/a_3411_1607# MAJ_0/a_644_83# UMA_1/a_3411_1607# MAJ_4/a_551_708# MAJ_5/w_26_1560#
+ MAJ_5/a_551_708# UMA_5/a_4705_1617# UMA_0/a_4705_1617# MAJ_3/a_1502_2030# MAJ_6/w_26_1560#
+ UMA_5/a_3411_1607# MAJ_6/a_551_708# UMA_0/a_3411_1607# MAJ_5/a_644_83# MAJ_1/a_644_83#
+ MAJ_7/w_26_1560# VSUBS
XMAJ_5 MAJ_5/w_26_1560# MAJ_5/a_551_708# UMA_5/a_n806_2017# m1_52380_205569# m1_52140_206158#
+ m1_52418_201623# MAJ_5/a_639_1698# UMA_5/a_3213_287# MAJ_5/a_644_83# m1_52180_202214#
+ UMA_5/a_121_287# MAJ_5/a_1502_2030# VSUBS MAJ_5/a_749_2028# MAJ
XMAJ_6 MAJ_6/w_26_1560# MAJ_6/a_551_708# UMA_6/a_n806_2017# m1_52379_209503# m1_52143_210093#
+ m1_52380_205569# MAJ_6/a_639_1698# UMA_6/a_3213_287# MAJ_6/a_644_83# m1_52140_206158#
+ UMA_6/a_121_287# MAJ_6/a_1502_2030# VSUBS MAJ_6/a_749_2028# MAJ
XMAJ_7 MAJ_7/w_26_1560# MAJ_7/a_551_708# UMA_7/a_n806_2017# MAJ_7/a_4594_2030# MAJ_7/a_3643_708#
+ m1_52379_209503# MAJ_7/a_639_1698# UMA_7/a_3213_287# MAJ_7/a_644_83# m1_52143_210093#
+ UMA_7/a_121_287# MAJ_7/a_1502_2030# VSUBS MAJ_7/a_749_2028# MAJ
XUMA_0 m1_53747_186215# UMA_0/a_4705_1617# UMA_0/a_209_1277# UMA_0/a_3411_1607# UMA_0/a_n806_2017#
+ UMA_0/a_n690_608# VSUBS UMA_0/a_121_287# UMA_0/m1_n6688_1443# m1_54160_186483# UMA_0/a_3213_287#
+ MAJ_0/w_26_1560# MAJ_0/a_749_2028# UMA_0/a_n912_608# UMA
XUMA_1 m1_53728_190208# UMA_1/a_4705_1617# UMA_1/a_209_1277# UMA_1/a_3411_1607# UMA_1/a_n806_2017#
+ m1_53747_186215# VSUBS UMA_1/a_121_287# m1_54160_186483# m1_54140_190478# UMA_1/a_3213_287#
+ MAJ_1/w_26_1560# MAJ_1/a_749_2028# UMA_1/a_n912_608# UMA
XUMA_2 m1_53670_194145# UMA_2/a_4705_1617# UMA_2/a_209_1277# UMA_2/a_3411_1607# UMA_2/a_n806_2017#
+ m1_53728_190208# VSUBS UMA_2/a_121_287# m1_54140_190478# m1_54085_194415# UMA_2/a_3213_287#
+ MAJ_2/w_26_1560# MAJ_2/a_749_2028# UMA_2/a_n912_608# UMA
XUMA_3 m1_53694_198104# UMA_3/a_4705_1617# UMA_3/a_209_1277# UMA_3/a_3411_1607# UMA_3/a_n806_2017#
+ m1_53670_194145# VSUBS UMA_3/a_121_287# m1_54085_194415# m1_54109_198374# UMA_3/a_3213_287#
+ MAJ_3/w_26_1560# MAJ_3/a_749_2028# UMA_3/a_n912_608# UMA
XUMA_5 m1_53690_205990# UMA_5/a_4705_1617# UMA_5/a_209_1277# UMA_5/a_3411_1607# UMA_5/a_n806_2017#
+ m1_53694_202051# VSUBS UMA_5/a_121_287# m1_54109_202321# m1_54107_206262# UMA_5/a_3213_287#
+ MAJ_5/w_26_1560# MAJ_5/a_749_2028# UMA_5/a_n912_608# UMA
XUMA_4 m1_53694_202051# UMA_4/a_4705_1617# UMA_4/a_209_1277# UMA_4/a_3411_1607# UMA_4/a_n806_2017#
+ m1_53694_198104# VSUBS UMA_4/a_121_287# m1_54109_198374# m1_54109_202321# UMA_4/a_3213_287#
+ MAJ_4/w_26_1560# MAJ_4/a_749_2028# UMA_4/a_n912_608# UMA
XUMA_6 m1_53630_209933# UMA_6/a_4705_1617# UMA_6/a_209_1277# UMA_6/a_3411_1607# UMA_6/a_n806_2017#
+ m1_53690_205990# VSUBS UMA_6/a_121_287# m1_54107_206262# m1_54045_210203# UMA_6/a_3213_287#
+ MAJ_6/w_26_1560# MAJ_6/a_749_2028# UMA_6/a_n912_608# UMA
XUMA_7 UMA_7/a_319_1607# UMA_7/a_4705_1617# UMA_7/a_209_1277# UMA_7/a_3411_1607# UMA_7/a_n806_2017#
+ m1_53630_209933# VSUBS UMA_7/a_121_287# m1_54045_210203# UMA_7/a_1613_1617# UMA_7/a_3213_287#
+ MAJ_7/w_26_1560# MAJ_7/a_749_2028# UMA_7/a_n912_608# UMA
XMAJ_0 MAJ_0/w_26_1560# MAJ_0/a_551_708# UMA_0/a_n806_2017# m1_52370_185794# m1_52134_186384#
+ MAJ_0/a_11429_1029# MAJ_0/a_639_1698# UMA_0/a_3213_287# MAJ_0/a_644_83# MAJ_0/m1_7413_2589#
+ UMA_0/a_121_287# MAJ_0/a_1502_2030# VSUBS MAJ_0/a_749_2028# MAJ
XMAJ_1 MAJ_1/w_26_1560# MAJ_1/a_551_708# UMA_1/a_n806_2017# m1_52370_189756# m1_52134_190346#
+ m1_52370_185794# MAJ_1/a_639_1698# UMA_1/a_3213_287# MAJ_1/a_644_83# m1_52134_186384#
+ UMA_1/a_121_287# MAJ_1/a_1502_2030# VSUBS MAJ_1/a_749_2028# MAJ
XMAJ_2 MAJ_2/w_26_1560# MAJ_2/a_551_708# UMA_2/a_n806_2017# m1_52351_193711# m1_52115_194301#
+ m1_52370_189756# MAJ_2/a_639_1698# UMA_2/a_3213_287# MAJ_2/a_644_83# m1_52134_190346#
+ UMA_2/a_121_287# MAJ_2/a_1502_2030# VSUBS MAJ_2/a_749_2028# MAJ
XMAJ_3 MAJ_3/w_26_1560# MAJ_3/a_551_708# UMA_3/a_n806_2017# m1_52410_197656# m1_52170_198245#
+ m1_52351_193711# MAJ_3/a_639_1698# UMA_3/a_3213_287# MAJ_3/a_644_83# m1_52115_194301#
+ UMA_3/a_121_287# MAJ_3/a_1502_2030# VSUBS MAJ_3/a_749_2028# MAJ
XMAJ_4 MAJ_4/w_26_1560# MAJ_4/a_551_708# UMA_4/a_n806_2017# m1_52418_201623# m1_52180_202214#
+ m1_52410_197656# MAJ_4/a_639_1698# UMA_4/a_3213_287# MAJ_4/a_644_83# m1_52170_198245#
+ UMA_4/a_121_287# MAJ_4/a_1502_2030# VSUBS MAJ_4/a_749_2028# MAJ
.ends

.subckt x16b_FA z z_not c0_b c0_not_b c15_not c15 s5_not s5 s0_not s0 s6_not s6 s1_not
+ s1 s7_not s7 s2_not s2 s8_not s8 s3_not s3 s9_not s9 s4_not s4 s10_not s10 s11_not
+ s11 s12_not s12 s13_not s13 s14_not s14 s15_not s15 c0_f c0_f_not vss vdd a0_f a0_not_f
+ b0 b0_not a1_f a1_not_f b1 b1_not a2_f a2_not_f b2 b2_not a3_f a3_not_f b3 b3_not
+ a4_f a4_not_f b4 b4_not a5_f a5_not_f b5 b5_not a6_f a6_not_f b6 b6_not a7_f a7_not_f
+ b7 b7_not a8_f a8_not_f b8 b8_not a9_f a9_not_f b9 b9_not a10_f a10_not_f b10 b10_not
+ a11_f a11_not_f b11 b11_not a12_f a12_not_f b12 b12_not a13_f a13_not_f b13 b13_not
+ a14_f a14_not_f b14 b14_not a15_f a15_not_f b15 b15_not a0_b a0_not_b a1_b a1_not_b
+ a2_b a2_not_b a3_b a3_not_b a4_b a4_not_b a5_b a5_not_b a6_b a6_not_b a7_b a7_not_b
+ a8_b a8_not_b a9_b a9_not_b a10_b a10_not_b a11_b a11_not_b a12_b a12_not_b a13_b
+ a13_not_b a14_b a14_not_b a15_b a15_not_b
X8b_FA_0 b8_not m1_12945_578# 8b_FA_0/UMA_4/a_4705_1617# b8 b13 8b_FA_0/UMA_4/a_3411_1607#
+ a_13565_n36782# a9_f a13_f a_13560_n35167# s12_not 8b_FA_0/MAJ_6/a_1502_2030# b14
+ a15_b m1_11125_463# a_13560_n35167# a14_b s12 a15_not_f a13_b vdd a14_not_f a12_b
+ a13_not_f a11_b b15_not a12_not_f 8b_FA_0/UMA_5/a_n912_608# a15_not_b a8_f a11_not_f
+ m1_11370_n128# a9_b vdd a14_not_b a10_not_f s8_not a8_b a12_f s13_not a9_not_f a13_not_b
+ b10 b14_not b15 a8_not_f m1_12525_313# a12_not_b s8 a11_not_b vdd s13 a10_not_b
+ a9_not_b b13_not a8_not_b vdd s9_not s14_not b12_not b11 a11_f vdd a_13565_n36782#
+ s9 a15_f s14 b11_not vdd b10_not s10_not s15_not b12 vdd 8b_FA_0/UMA_5/a_3411_1607#
+ 8b_FA_0/MAJ_6/a_551_708# s15 a10_f 8b_FA_0/MAJ_1/a_644_83# vdd vss x8b_FA
X8b_FA_1 b0_not c0_not_b s3_not b0 b5 s3 m1_12525_313# a1_f a5_f m1_12945_578# s4_not
+ b1 b6 a7_b 8b_FA_1/MAJ_7/a_3643_708# m1_11125_463# a6_b 8b_FA_1/UMA_3/a_3411_1607#
+ a7_not_f a5_b vdd a6_not_f a4_b a5_not_f a3_b b7_not a4_not_f a2_b a7_not_b a0_f
+ a3_not_f c0_f a1_b vdd a6_not_b a2_not_f 8b_FA_1/UMA_7/a_4705_1617# a0_b a4_f 8b_FA_1/UMA_2/a_4705_1617#
+ a1_not_f a5_not_b b2 b6_not b7 a0_not_f c0_b a4_not_b 8b_FA_1/UMA_7/a_3411_1607#
+ a3_not_b vdd 8b_FA_1/UMA_2/a_3411_1607# a2_not_b a1_not_b b5_not a0_not_b vdd s1_not
+ s6_not 8b_FA_1/MAJ_3/a_551_708# b3 8b_FA_1/MAJ_4/a_644_83# vdd m1_11370_n128# s1
+ a7_f s6 b3_not vdd b2_not s2_not s7_not b4 vdd s2 b1_not s7 a2_f a6_f vdd vss x8b_FA
X0 z a_13560_n35167# c15 vss nfet_03v3 ad=0.65797p pd=3.76u as=0.74287p ps=3.88u w=1.415u l=0.55u
X1 c15 a_13560_n35167# z_not vdd pfet_03v3 ad=0.6669p pd=3.55u as=0.60515p ps=3.45u w=1.235u l=0.5u
X2 z_not a_13565_n36782# c15_not vdd pfet_03v3 ad=0.70395p pd=3.61u as=0.6422p ps=3.51u w=1.235u l=0.5u
X3 c15_not a_13565_n36782# z vss nfet_03v3 ad=0.64155p pd=3.67u as=0.64837p ps=3.68u w=1.365u l=0.55u
X4 z_not a_13560_n35167# c15_not vss nfet_03v3 ad=0.6925p pd=3.77u as=0.67172p ps=3.74u w=1.385u l=0.55u
X5 z a_13565_n36782# c15 vdd pfet_03v3 ad=0.60515p pd=3.45u as=0.6669p ps=3.55u w=1.235u l=0.5u
X6 c15 a_13565_n36782# z_not vss nfet_03v3 ad=0.6576p pd=3.7u as=0.63705p ps=3.67u w=1.37u l=0.55u
X7 c15_not a_13560_n35167# z vdd pfet_03v3 ad=0.60515p pd=3.45u as=0.64837p ps=3.52u w=1.235u l=0.5u
.ends

