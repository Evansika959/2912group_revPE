VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fa8b_rev
  CLASS BLOCK ;
  FOREIGN fa8b_rev ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.665 BY 212.100 ;
  PIN c_8_not
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 104.010 24.915 108.095 25.250 ;
    END
  END c_8_not
  PIN z
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 100.280 27.290 111.325 27.590 ;
    END
  END z
  PIN z_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT 102.630 26.755 108.680 27.025 ;
    END
  END z_not
  PIN c0
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 161.170 184.800 164.390 185.100 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 30.005 181.695 50.350 181.990 ;
    END
  END c0
  PIN c0_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 158.225 184.055 165.950 184.355 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 29.825 180.830 50.935 181.125 ;
    END
  END c0_not
  PIN s0
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 152.405 180.965 162.485 181.300 ;
    END
  END s0
  PIN s0_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 159.755 183.040 162.485 183.315 ;
    END
  END s0_not
  PIN s1
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 152.205 161.240 162.285 161.575 ;
    END
  END s1
  PIN s1_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 159.555 163.315 162.285 163.590 ;
    END
  END s1_not
  PIN s2
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 152.360 141.595 162.440 141.930 ;
    END
  END s2
  PIN s2_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 159.710 143.670 162.440 143.945 ;
    END
  END s2_not
  PIN s3
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 152.360 121.800 162.440 122.135 ;
    END
  END s3
  PIN s3_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 159.710 123.875 162.440 124.150 ;
    END
  END s3_not
  PIN s4
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 152.280 102.045 162.360 102.380 ;
    END
  END s4
  PIN s4_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 159.630 104.120 162.360 104.395 ;
    END
  END s4_not
  PIN s5
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 152.385 82.330 162.465 82.665 ;
    END
  END s5
  PIN s5_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 159.735 84.405 162.465 84.680 ;
    END
  END s5_not
  PIN s6
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 152.385 62.360 162.465 62.695 ;
    END
  END s6
  PIN s6_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 159.735 64.435 162.465 64.710 ;
    END
  END s6_not
  PIN s7
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 152.385 42.695 162.465 43.030 ;
    END
  END s7
  PIN s7_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 159.735 44.770 162.465 45.045 ;
    END
  END s7_not
  PIN c_8
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal3 ;
        RECT 118.430 18.370 119.455 18.720 ;
    END
  END c_8
  PIN a0_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 32.960 184.850 35.420 185.155 ;
    END
  END a0_f
  PIN a0_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 32.920 184.115 35.425 184.410 ;
    END
  END a0_not_f
  PIN a0_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 146.970 189.670 162.705 190.080 ;
    END
  END a0_b
  PIN a0_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 147.565 188.890 162.695 189.345 ;
    END
  END a0_not_b
  PIN a7_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 32.830 46.535 35.290 46.840 ;
    END
  END a7_f
  PIN a7_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 32.790 45.800 35.295 46.095 ;
    END
  END a7_not_f
  PIN a7_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 146.950 51.400 162.685 51.810 ;
    END
  END a7_b
  PIN a7_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 147.545 50.620 162.675 51.075 ;
    END
  END a7_not_b
  PIN b0
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 32.925 183.400 35.440 183.695 ;
    END
  END b0
  PIN b0_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 32.960 182.770 35.425 183.065 ;
    END
  END b0_not
  PIN a1
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 32.915 165.160 35.375 165.465 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 146.770 169.945 162.505 170.355 ;
    END
  END a1
  PIN a1_not
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 32.875 164.425 35.380 164.720 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 147.365 169.165 162.495 169.620 ;
    END
  END a1_not
  PIN b1
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 32.880 163.710 35.395 164.005 ;
    END
  END b1
  PIN b1_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 32.915 163.080 35.380 163.375 ;
    END
  END b1_not
  PIN a2
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 33.105 145.450 35.565 145.755 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 146.925 150.300 162.660 150.710 ;
    END
  END a2
  PIN a2_not
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 33.065 144.715 35.570 145.010 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 147.520 149.520 162.650 149.975 ;
    END
  END a2_not
  PIN b2
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 33.070 144.000 35.585 144.295 ;
    END
  END b2
  PIN b2_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 33.105 143.370 35.570 143.665 ;
    END
  END b2_not
  PIN a3
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 32.910 125.610 35.370 125.915 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 146.925 130.505 162.660 130.915 ;
    END
  END a3
  PIN a3_not
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 32.870 124.875 35.375 125.170 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 147.520 129.725 162.650 130.180 ;
    END
  END a3_not
  PIN b3
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 32.875 124.160 35.390 124.455 ;
    END
  END b3
  PIN b3_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 32.910 123.530 35.375 123.825 ;
    END
  END b3_not
  PIN a4
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 32.780 105.900 35.240 106.205 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 146.845 110.750 162.580 111.160 ;
    END
  END a4
  PIN a4_not
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 32.740 105.165 35.245 105.460 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 147.440 109.970 162.570 110.425 ;
    END
  END a4_not
  PIN b4
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 32.745 104.450 35.260 104.745 ;
    END
  END b4
  PIN b4_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 32.780 103.820 35.245 104.115 ;
    END
  END b4_not
  PIN a5
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 32.910 86.140 35.370 86.445 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 146.950 91.035 162.685 91.445 ;
    END
  END a5
  PIN a5_not
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 32.870 85.405 35.375 85.700 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 147.545 90.255 162.675 90.710 ;
    END
  END a5_not
  PIN b5
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 32.875 84.690 35.390 84.985 ;
    END
  END b5
  PIN b5_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 32.910 84.060 35.375 84.355 ;
    END
  END b5_not
  PIN a6
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 32.860 66.330 35.320 66.635 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 146.950 71.065 162.685 71.475 ;
    END
  END a6
  PIN a6_not
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 32.820 65.595 35.325 65.890 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 147.545 70.285 162.675 70.740 ;
    END
  END a6_not
  PIN b6
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 32.825 64.880 35.340 65.175 ;
    END
  END b6
  PIN b6_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 32.860 64.250 35.325 64.545 ;
    END
  END b6_not
  PIN b7
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 32.795 45.085 35.310 45.380 ;
    END
  END b7
  PIN b7_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 32.830 44.455 35.295 44.750 ;
    END
  END b7_not
  OBS
      LAYER Nwell ;
        RECT 33.240 19.365 162.485 191.395 ;
      LAYER Metal1 ;
        RECT 33.670 185.400 170.510 191.395 ;
        RECT 33.670 184.655 160.870 185.400 ;
        RECT 164.690 184.655 170.510 185.400 ;
        RECT 33.670 183.755 157.925 184.655 ;
        RECT 166.250 183.755 170.510 184.655 ;
        RECT 33.670 183.615 170.510 183.755 ;
        RECT 33.670 182.740 159.455 183.615 ;
        RECT 162.785 182.740 170.510 183.615 ;
        RECT 33.670 181.600 170.510 182.740 ;
        RECT 33.670 180.665 152.105 181.600 ;
        RECT 162.785 180.665 170.510 181.600 ;
        RECT 33.670 163.890 170.510 180.665 ;
        RECT 33.670 163.015 159.255 163.890 ;
        RECT 162.585 163.015 170.510 163.890 ;
        RECT 33.670 161.875 170.510 163.015 ;
        RECT 33.670 160.940 151.905 161.875 ;
        RECT 162.585 160.940 170.510 161.875 ;
        RECT 33.670 144.245 170.510 160.940 ;
        RECT 33.670 143.370 159.410 144.245 ;
        RECT 162.740 143.370 170.510 144.245 ;
        RECT 33.670 142.230 170.510 143.370 ;
        RECT 33.670 141.295 152.060 142.230 ;
        RECT 162.740 141.295 170.510 142.230 ;
        RECT 33.670 124.450 170.510 141.295 ;
        RECT 33.670 123.575 159.410 124.450 ;
        RECT 162.740 123.575 170.510 124.450 ;
        RECT 33.670 122.435 170.510 123.575 ;
        RECT 33.670 121.500 152.060 122.435 ;
        RECT 162.740 121.500 170.510 122.435 ;
        RECT 33.670 104.695 170.510 121.500 ;
        RECT 33.670 103.820 159.330 104.695 ;
        RECT 162.660 103.820 170.510 104.695 ;
        RECT 33.670 102.680 170.510 103.820 ;
        RECT 33.670 101.745 151.980 102.680 ;
        RECT 162.660 101.745 170.510 102.680 ;
        RECT 33.670 84.980 170.510 101.745 ;
        RECT 33.670 84.105 159.435 84.980 ;
        RECT 162.765 84.105 170.510 84.980 ;
        RECT 33.670 82.965 170.510 84.105 ;
        RECT 33.670 82.030 152.085 82.965 ;
        RECT 162.765 82.030 170.510 82.965 ;
        RECT 33.670 65.010 170.510 82.030 ;
        RECT 33.670 64.135 159.435 65.010 ;
        RECT 162.765 64.135 170.510 65.010 ;
        RECT 33.670 62.995 170.510 64.135 ;
        RECT 33.670 62.060 152.085 62.995 ;
        RECT 162.765 62.060 170.510 62.995 ;
        RECT 33.670 45.345 170.510 62.060 ;
        RECT 33.670 44.470 159.435 45.345 ;
        RECT 162.765 44.470 170.510 45.345 ;
        RECT 33.670 43.330 170.510 44.470 ;
        RECT 33.670 42.395 152.085 43.330 ;
        RECT 162.765 42.395 170.510 43.330 ;
        RECT 33.670 27.890 170.510 42.395 ;
        RECT 33.670 26.990 99.980 27.890 ;
        RECT 111.625 26.990 170.510 27.890 ;
        RECT 33.670 26.455 102.330 26.990 ;
        RECT 108.980 26.455 170.510 26.990 ;
        RECT 33.670 25.550 170.510 26.455 ;
        RECT 33.670 24.615 103.710 25.550 ;
        RECT 108.395 24.615 170.510 25.550 ;
        RECT 33.670 19.360 170.510 24.615 ;
      LAYER Metal2 ;
        RECT 29.910 7.790 165.840 191.395 ;
      LAYER Metal3 ;
        RECT 12.415 190.380 181.500 204.855 ;
        RECT 12.415 189.370 146.670 190.380 ;
        RECT 163.005 189.370 181.500 190.380 ;
        RECT 12.415 188.590 147.265 189.370 ;
        RECT 162.995 188.590 181.500 189.370 ;
        RECT 12.415 185.455 181.500 188.590 ;
        RECT 12.415 184.710 32.660 185.455 ;
        RECT 35.720 184.710 181.500 185.455 ;
        RECT 12.415 183.815 32.620 184.710 ;
        RECT 35.725 183.995 181.500 184.710 ;
        RECT 12.415 183.100 32.625 183.815 ;
        RECT 35.740 183.100 181.500 183.995 ;
        RECT 12.415 182.470 32.660 183.100 ;
        RECT 35.725 182.470 181.500 183.100 ;
        RECT 12.415 182.290 181.500 182.470 ;
        RECT 12.415 181.425 29.705 182.290 ;
        RECT 50.650 181.425 181.500 182.290 ;
        RECT 12.415 180.530 29.525 181.425 ;
        RECT 51.235 180.530 181.500 181.425 ;
        RECT 12.415 170.655 181.500 180.530 ;
        RECT 12.415 169.645 146.470 170.655 ;
        RECT 162.805 169.645 181.500 170.655 ;
        RECT 12.415 168.865 147.065 169.645 ;
        RECT 162.795 168.865 181.500 169.645 ;
        RECT 12.415 165.765 181.500 168.865 ;
        RECT 12.415 165.020 32.615 165.765 ;
        RECT 35.675 165.020 181.500 165.765 ;
        RECT 12.415 164.125 32.575 165.020 ;
        RECT 35.680 164.305 181.500 165.020 ;
        RECT 12.415 163.410 32.580 164.125 ;
        RECT 35.695 163.410 181.500 164.305 ;
        RECT 12.415 162.780 32.615 163.410 ;
        RECT 35.680 162.780 181.500 163.410 ;
        RECT 12.415 151.010 181.500 162.780 ;
        RECT 12.415 150.000 146.625 151.010 ;
        RECT 162.960 150.000 181.500 151.010 ;
        RECT 12.415 149.220 147.220 150.000 ;
        RECT 162.950 149.220 181.500 150.000 ;
        RECT 12.415 146.055 181.500 149.220 ;
        RECT 12.415 145.310 32.805 146.055 ;
        RECT 35.865 145.310 181.500 146.055 ;
        RECT 12.415 144.415 32.765 145.310 ;
        RECT 35.870 144.595 181.500 145.310 ;
        RECT 12.415 143.700 32.770 144.415 ;
        RECT 35.885 143.700 181.500 144.595 ;
        RECT 12.415 143.070 32.805 143.700 ;
        RECT 35.870 143.070 181.500 143.700 ;
        RECT 12.415 131.215 181.500 143.070 ;
        RECT 12.415 130.205 146.625 131.215 ;
        RECT 162.960 130.205 181.500 131.215 ;
        RECT 12.415 129.425 147.220 130.205 ;
        RECT 162.950 129.425 181.500 130.205 ;
        RECT 12.415 126.215 181.500 129.425 ;
        RECT 12.415 125.470 32.610 126.215 ;
        RECT 35.670 125.470 181.500 126.215 ;
        RECT 12.415 124.575 32.570 125.470 ;
        RECT 35.675 124.755 181.500 125.470 ;
        RECT 12.415 123.860 32.575 124.575 ;
        RECT 35.690 123.860 181.500 124.755 ;
        RECT 12.415 123.230 32.610 123.860 ;
        RECT 35.675 123.230 181.500 123.860 ;
        RECT 12.415 111.460 181.500 123.230 ;
        RECT 12.415 110.450 146.545 111.460 ;
        RECT 162.880 110.450 181.500 111.460 ;
        RECT 12.415 109.670 147.140 110.450 ;
        RECT 162.870 109.670 181.500 110.450 ;
        RECT 12.415 106.505 181.500 109.670 ;
        RECT 12.415 105.760 32.480 106.505 ;
        RECT 35.540 105.760 181.500 106.505 ;
        RECT 12.415 104.865 32.440 105.760 ;
        RECT 35.545 105.045 181.500 105.760 ;
        RECT 12.415 104.150 32.445 104.865 ;
        RECT 35.560 104.150 181.500 105.045 ;
        RECT 12.415 103.520 32.480 104.150 ;
        RECT 35.545 103.520 181.500 104.150 ;
        RECT 12.415 91.745 181.500 103.520 ;
        RECT 12.415 90.735 146.650 91.745 ;
        RECT 162.985 90.735 181.500 91.745 ;
        RECT 12.415 89.955 147.245 90.735 ;
        RECT 162.975 89.955 181.500 90.735 ;
        RECT 12.415 86.745 181.500 89.955 ;
        RECT 12.415 86.000 32.610 86.745 ;
        RECT 35.670 86.000 181.500 86.745 ;
        RECT 12.415 85.105 32.570 86.000 ;
        RECT 35.675 85.285 181.500 86.000 ;
        RECT 12.415 84.390 32.575 85.105 ;
        RECT 35.690 84.390 181.500 85.285 ;
        RECT 12.415 83.760 32.610 84.390 ;
        RECT 35.675 83.760 181.500 84.390 ;
        RECT 12.415 71.775 181.500 83.760 ;
        RECT 12.415 70.765 146.650 71.775 ;
        RECT 162.985 70.765 181.500 71.775 ;
        RECT 12.415 69.985 147.245 70.765 ;
        RECT 162.975 69.985 181.500 70.765 ;
        RECT 12.415 66.935 181.500 69.985 ;
        RECT 12.415 66.190 32.560 66.935 ;
        RECT 35.620 66.190 181.500 66.935 ;
        RECT 12.415 65.295 32.520 66.190 ;
        RECT 35.625 65.475 181.500 66.190 ;
        RECT 12.415 64.580 32.525 65.295 ;
        RECT 35.640 64.580 181.500 65.475 ;
        RECT 12.415 63.950 32.560 64.580 ;
        RECT 35.625 63.950 181.500 64.580 ;
        RECT 12.415 52.110 181.500 63.950 ;
        RECT 12.415 51.100 146.650 52.110 ;
        RECT 162.985 51.100 181.500 52.110 ;
        RECT 12.415 50.320 147.245 51.100 ;
        RECT 162.975 50.320 181.500 51.100 ;
        RECT 12.415 47.140 181.500 50.320 ;
        RECT 12.415 46.395 32.530 47.140 ;
        RECT 35.590 46.395 181.500 47.140 ;
        RECT 12.415 45.500 32.490 46.395 ;
        RECT 35.595 45.680 181.500 46.395 ;
        RECT 12.415 44.785 32.495 45.500 ;
        RECT 35.610 44.785 181.500 45.680 ;
        RECT 12.415 44.155 32.530 44.785 ;
        RECT 35.595 44.155 181.500 44.785 ;
        RECT 12.415 19.020 181.500 44.155 ;
        RECT 12.415 18.070 118.130 19.020 ;
        RECT 119.755 18.070 181.500 19.020 ;
        RECT 12.415 7.790 181.500 18.070 ;
      LAYER Metal4 ;
        RECT 17.210 7.745 180.600 204.920 ;
  END
END fa8b_rev
END LIBRARY

